-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_727_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_723_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_1 : boolean;
  signal type_cast_1280_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1060_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_741_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1396_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1010_inst_req_1 : boolean;
  signal if_stmt_632_branch_ack_1 : boolean;
  signal type_cast_727_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1390_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1010_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 : boolean;
  signal addr_of_689_final_reg_ack_1 : boolean;
  signal type_cast_592_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_ack_0 : boolean;
  signal type_cast_592_inst_req_0 : boolean;
  signal type_cast_538_inst_ack_1 : boolean;
  signal type_cast_538_inst_req_1 : boolean;
  signal type_cast_538_inst_ack_0 : boolean;
  signal type_cast_538_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_ack_1 : boolean;
  signal type_cast_709_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_588_inst_req_0 : boolean;
  signal type_cast_38_inst_req_0 : boolean;
  signal type_cast_38_inst_ack_0 : boolean;
  signal type_cast_38_inst_req_1 : boolean;
  signal type_cast_38_inst_ack_1 : boolean;
  signal type_cast_709_inst_req_1 : boolean;
  signal type_cast_727_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_1 : boolean;
  signal type_cast_1048_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 : boolean;
  signal addr_of_689_final_reg_req_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_1 : boolean;
  signal type_cast_610_inst_ack_0 : boolean;
  signal type_cast_1328_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 : boolean;
  signal addr_of_689_final_reg_req_1 : boolean;
  signal WPIPE_Block1_start_1016_inst_req_1 : boolean;
  signal type_cast_51_inst_req_0 : boolean;
  signal type_cast_51_inst_ack_0 : boolean;
  signal type_cast_51_inst_req_1 : boolean;
  signal type_cast_51_inst_ack_1 : boolean;
  signal type_cast_727_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_705_inst_req_0 : boolean;
  signal type_cast_63_inst_req_0 : boolean;
  signal type_cast_63_inst_ack_0 : boolean;
  signal type_cast_63_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_1 : boolean;
  signal ptr_deref_618_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 : boolean;
  signal if_stmt_632_branch_req_0 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal array_obj_ref_688_index_offset_ack_1 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal ptr_deref_618_store_0_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_0 : boolean;
  signal WPIPE_Block0_start_990_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_692_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 : boolean;
  signal type_cast_610_inst_ack_1 : boolean;
  signal type_cast_88_inst_req_0 : boolean;
  signal type_cast_88_inst_ack_0 : boolean;
  signal array_obj_ref_688_index_offset_req_1 : boolean;
  signal type_cast_88_inst_req_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_0 : boolean;
  signal type_cast_88_inst_ack_1 : boolean;
  signal type_cast_709_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1069_inst_ack_1 : boolean;
  signal addr_of_1310_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 : boolean;
  signal type_cast_659_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_req_0 : boolean;
  signal type_cast_610_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1010_inst_ack_1 : boolean;
  signal type_cast_101_inst_req_0 : boolean;
  signal WPIPE_Block0_start_984_inst_req_0 : boolean;
  signal type_cast_101_inst_ack_0 : boolean;
  signal type_cast_101_inst_req_1 : boolean;
  signal type_cast_101_inst_ack_1 : boolean;
  signal type_cast_709_inst_req_0 : boolean;
  signal type_cast_574_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_996_inst_req_1 : boolean;
  signal type_cast_659_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 : boolean;
  signal type_cast_574_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 : boolean;
  signal addr_of_689_final_reg_ack_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_ack_1 : boolean;
  signal type_cast_113_inst_req_0 : boolean;
  signal type_cast_113_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_1 : boolean;
  signal ptr_deref_618_store_0_ack_0 : boolean;
  signal type_cast_113_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_1 : boolean;
  signal ptr_deref_618_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_req_0 : boolean;
  signal array_obj_ref_688_index_offset_ack_0 : boolean;
  signal type_cast_126_inst_req_0 : boolean;
  signal type_cast_126_inst_ack_0 : boolean;
  signal type_cast_659_inst_ack_0 : boolean;
  signal type_cast_126_inst_req_1 : boolean;
  signal type_cast_126_inst_ack_1 : boolean;
  signal type_cast_574_inst_ack_0 : boolean;
  signal type_cast_659_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 : boolean;
  signal type_cast_339_inst_req_0 : boolean;
  signal type_cast_339_inst_ack_0 : boolean;
  signal type_cast_339_inst_req_1 : boolean;
  signal type_cast_339_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_348_inst_ack_1 : boolean;
  signal type_cast_138_inst_req_0 : boolean;
  signal type_cast_138_inst_ack_0 : boolean;
  signal type_cast_138_inst_req_1 : boolean;
  signal type_cast_138_inst_ack_1 : boolean;
  signal type_cast_574_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1057_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 : boolean;
  signal type_cast_696_inst_ack_1 : boolean;
  signal type_cast_696_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_ack_0 : boolean;
  signal type_cast_610_inst_req_0 : boolean;
  signal array_obj_ref_688_index_offset_req_0 : boolean;
  signal type_cast_151_inst_req_0 : boolean;
  signal type_cast_151_inst_ack_0 : boolean;
  signal type_cast_151_inst_req_1 : boolean;
  signal type_cast_151_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_1 : boolean;
  signal type_cast_163_inst_req_0 : boolean;
  signal type_cast_163_inst_ack_0 : boolean;
  signal type_cast_163_inst_req_1 : boolean;
  signal type_cast_1048_inst_ack_0 : boolean;
  signal type_cast_163_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_972_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 : boolean;
  signal type_cast_696_inst_ack_0 : boolean;
  signal type_cast_696_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1013_inst_ack_0 : boolean;
  signal type_cast_176_inst_req_0 : boolean;
  signal type_cast_176_inst_ack_0 : boolean;
  signal type_cast_176_inst_req_1 : boolean;
  signal type_cast_176_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1396_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 : boolean;
  signal type_cast_1328_inst_req_0 : boolean;
  signal type_cast_188_inst_req_0 : boolean;
  signal type_cast_188_inst_ack_0 : boolean;
  signal type_cast_188_inst_req_1 : boolean;
  signal type_cast_188_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1057_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_0 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_972_inst_req_1 : boolean;
  signal type_cast_201_inst_req_0 : boolean;
  signal type_cast_201_inst_ack_0 : boolean;
  signal type_cast_201_inst_req_1 : boolean;
  signal type_cast_201_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_570_inst_req_0 : boolean;
  signal WPIPE_Block0_start_975_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1057_inst_req_1 : boolean;
  signal type_cast_210_inst_req_0 : boolean;
  signal type_cast_210_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_req_1 : boolean;
  signal type_cast_210_inst_req_1 : boolean;
  signal type_cast_210_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1000_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1013_inst_req_1 : boolean;
  signal type_cast_214_inst_req_0 : boolean;
  signal type_cast_214_inst_ack_0 : boolean;
  signal type_cast_214_inst_req_1 : boolean;
  signal type_cast_214_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_req_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_1 : boolean;
  signal type_cast_218_inst_req_0 : boolean;
  signal type_cast_218_inst_ack_0 : boolean;
  signal type_cast_218_inst_req_1 : boolean;
  signal type_cast_218_inst_ack_1 : boolean;
  signal type_cast_556_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_req_1 : boolean;
  signal type_cast_1048_inst_req_1 : boolean;
  signal type_cast_255_inst_req_0 : boolean;
  signal type_cast_255_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_ack_0 : boolean;
  signal type_cast_255_inst_req_1 : boolean;
  signal type_cast_255_inst_ack_1 : boolean;
  signal type_cast_556_inst_req_1 : boolean;
  signal type_cast_259_inst_req_0 : boolean;
  signal type_cast_259_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_534_inst_req_0 : boolean;
  signal type_cast_259_inst_req_1 : boolean;
  signal type_cast_259_inst_ack_1 : boolean;
  signal type_cast_556_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_606_inst_req_0 : boolean;
  signal type_cast_263_inst_req_0 : boolean;
  signal type_cast_263_inst_ack_0 : boolean;
  signal type_cast_263_inst_req_1 : boolean;
  signal type_cast_263_inst_ack_1 : boolean;
  signal type_cast_556_inst_req_0 : boolean;
  signal type_cast_267_inst_req_0 : boolean;
  signal type_cast_1048_inst_ack_1 : boolean;
  signal type_cast_267_inst_ack_0 : boolean;
  signal type_cast_267_inst_req_1 : boolean;
  signal type_cast_267_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_996_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_285_inst_ack_1 : boolean;
  signal type_cast_289_inst_req_0 : boolean;
  signal type_cast_289_inst_ack_0 : boolean;
  signal type_cast_289_inst_req_1 : boolean;
  signal type_cast_289_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_298_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1057_inst_ack_1 : boolean;
  signal type_cast_302_inst_req_0 : boolean;
  signal type_cast_302_inst_ack_0 : boolean;
  signal type_cast_302_inst_req_1 : boolean;
  signal type_cast_302_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_310_inst_ack_1 : boolean;
  signal type_cast_1378_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1013_inst_ack_1 : boolean;
  signal type_cast_592_inst_ack_1 : boolean;
  signal type_cast_592_inst_req_1 : boolean;
  signal type_cast_314_inst_req_0 : boolean;
  signal type_cast_314_inst_ack_0 : boolean;
  signal type_cast_314_inst_req_1 : boolean;
  signal type_cast_314_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_552_inst_req_0 : boolean;
  signal if_stmt_632_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_323_inst_ack_1 : boolean;
  signal type_cast_327_inst_req_0 : boolean;
  signal type_cast_327_inst_ack_0 : boolean;
  signal type_cast_327_inst_req_1 : boolean;
  signal type_cast_327_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_975_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_335_inst_ack_1 : boolean;
  signal type_cast_352_inst_req_0 : boolean;
  signal type_cast_352_inst_ack_0 : boolean;
  signal type_cast_352_inst_req_1 : boolean;
  signal type_cast_352_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_360_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_984_inst_req_1 : boolean;
  signal type_cast_364_inst_req_0 : boolean;
  signal type_cast_364_inst_ack_0 : boolean;
  signal type_cast_364_inst_req_1 : boolean;
  signal type_cast_364_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1050_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_373_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1050_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_1 : boolean;
  signal type_cast_377_inst_req_0 : boolean;
  signal type_cast_377_inst_ack_0 : boolean;
  signal type_cast_377_inst_req_1 : boolean;
  signal type_cast_377_inst_ack_1 : boolean;
  signal addr_of_1310_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1050_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_385_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_0 : boolean;
  signal type_cast_389_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1050_inst_ack_1 : boolean;
  signal type_cast_389_inst_ack_0 : boolean;
  signal type_cast_389_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1016_inst_req_0 : boolean;
  signal type_cast_389_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_398_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_req_0 : boolean;
  signal type_cast_402_inst_req_0 : boolean;
  signal type_cast_402_inst_ack_0 : boolean;
  signal addr_of_1310_final_reg_ack_1 : boolean;
  signal type_cast_402_inst_req_1 : boolean;
  signal type_cast_402_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1016_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_993_inst_req_1 : boolean;
  signal WPIPE_Block0_start_978_inst_req_1 : boolean;
  signal if_stmt_416_branch_req_0 : boolean;
  signal if_stmt_416_branch_ack_1 : boolean;
  signal if_stmt_416_branch_ack_0 : boolean;
  signal if_stmt_431_branch_req_0 : boolean;
  signal if_stmt_431_branch_ack_1 : boolean;
  signal if_stmt_431_branch_ack_0 : boolean;
  signal type_cast_452_inst_req_0 : boolean;
  signal type_cast_452_inst_ack_0 : boolean;
  signal type_cast_452_inst_req_1 : boolean;
  signal type_cast_452_inst_ack_1 : boolean;
  signal array_obj_ref_481_index_offset_req_0 : boolean;
  signal array_obj_ref_481_index_offset_ack_0 : boolean;
  signal array_obj_ref_481_index_offset_req_1 : boolean;
  signal array_obj_ref_481_index_offset_ack_1 : boolean;
  signal addr_of_482_final_reg_req_0 : boolean;
  signal addr_of_482_final_reg_ack_0 : boolean;
  signal addr_of_482_final_reg_req_1 : boolean;
  signal addr_of_482_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_485_inst_ack_1 : boolean;
  signal type_cast_489_inst_req_0 : boolean;
  signal type_cast_489_inst_ack_0 : boolean;
  signal type_cast_489_inst_req_1 : boolean;
  signal type_cast_489_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_498_inst_ack_1 : boolean;
  signal type_cast_502_inst_req_0 : boolean;
  signal type_cast_502_inst_ack_0 : boolean;
  signal type_cast_502_inst_req_1 : boolean;
  signal type_cast_502_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_516_inst_ack_1 : boolean;
  signal type_cast_520_inst_req_0 : boolean;
  signal type_cast_520_inst_ack_0 : boolean;
  signal type_cast_520_inst_req_1 : boolean;
  signal type_cast_520_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1060_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1069_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_ack_1 : boolean;
  signal type_cast_745_inst_req_0 : boolean;
  signal type_cast_745_inst_ack_0 : boolean;
  signal type_cast_745_inst_req_1 : boolean;
  signal type_cast_745_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_759_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1393_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1010_inst_req_0 : boolean;
  signal type_cast_763_inst_req_0 : boolean;
  signal type_cast_763_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1066_inst_req_1 : boolean;
  signal type_cast_763_inst_req_1 : boolean;
  signal type_cast_763_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1399_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1396_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1060_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1034_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1034_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_777_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1069_inst_ack_0 : boolean;
  signal type_cast_781_inst_req_0 : boolean;
  signal type_cast_781_inst_ack_0 : boolean;
  signal type_cast_781_inst_req_1 : boolean;
  signal type_cast_781_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1060_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1034_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1034_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_795_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1393_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1069_inst_req_0 : boolean;
  signal type_cast_799_inst_req_0 : boolean;
  signal type_cast_799_inst_ack_0 : boolean;
  signal type_cast_799_inst_req_1 : boolean;
  signal type_cast_799_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_813_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1007_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_ack_0 : boolean;
  signal type_cast_817_inst_req_0 : boolean;
  signal type_cast_817_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1066_inst_req_0 : boolean;
  signal type_cast_817_inst_req_1 : boolean;
  signal type_cast_817_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_ack_1 : boolean;
  signal type_cast_1055_inst_ack_1 : boolean;
  signal type_cast_1055_inst_req_1 : boolean;
  signal type_cast_1280_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1007_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_1 : boolean;
  signal WPIPE_Block0_start_996_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_996_inst_req_0 : boolean;
  signal ptr_deref_825_store_0_req_0 : boolean;
  signal WPIPE_Block0_start_1007_inst_ack_0 : boolean;
  signal ptr_deref_825_store_0_ack_0 : boolean;
  signal ptr_deref_825_store_0_req_1 : boolean;
  signal WPIPE_Block0_start_1007_inst_req_0 : boolean;
  signal ptr_deref_825_store_0_ack_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_ack_1 : boolean;
  signal if_stmt_839_branch_req_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_1 : boolean;
  signal if_stmt_839_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_0 : boolean;
  signal WPIPE_Block0_start_981_inst_req_1 : boolean;
  signal if_stmt_839_branch_ack_0 : boolean;
  signal type_cast_850_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_0 : boolean;
  signal type_cast_850_inst_ack_0 : boolean;
  signal type_cast_850_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_0 : boolean;
  signal type_cast_850_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_req_1 : boolean;
  signal type_cast_854_inst_req_0 : boolean;
  signal type_cast_854_inst_ack_0 : boolean;
  signal type_cast_1328_inst_req_1 : boolean;
  signal type_cast_854_inst_req_1 : boolean;
  signal type_cast_854_inst_ack_1 : boolean;
  signal type_cast_1378_inst_req_0 : boolean;
  signal type_cast_1055_inst_ack_0 : boolean;
  signal type_cast_1280_inst_ack_1 : boolean;
  signal type_cast_1055_inst_req_0 : boolean;
  signal type_cast_858_inst_req_0 : boolean;
  signal type_cast_858_inst_ack_0 : boolean;
  signal type_cast_858_inst_req_1 : boolean;
  signal type_cast_858_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1402_inst_req_0 : boolean;
  signal if_stmt_876_branch_req_0 : boolean;
  signal WPIPE_Block0_start_1004_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_0 : boolean;
  signal if_stmt_876_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_req_0 : boolean;
  signal if_stmt_876_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_1 : boolean;
  signal type_cast_903_inst_req_0 : boolean;
  signal type_cast_903_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1402_inst_ack_0 : boolean;
  signal type_cast_903_inst_req_1 : boolean;
  signal type_cast_903_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1072_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1004_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1004_inst_ack_0 : boolean;
  signal array_obj_ref_932_index_offset_req_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_1 : boolean;
  signal array_obj_ref_932_index_offset_ack_0 : boolean;
  signal array_obj_ref_932_index_offset_req_1 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_1 : boolean;
  signal array_obj_ref_932_index_offset_ack_1 : boolean;
  signal WPIPE_Block0_start_1004_inst_req_0 : boolean;
  signal addr_of_933_final_reg_req_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_0 : boolean;
  signal addr_of_933_final_reg_ack_0 : boolean;
  signal addr_of_933_final_reg_req_1 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_0 : boolean;
  signal addr_of_933_final_reg_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_0 : boolean;
  signal ptr_deref_936_store_0_req_0 : boolean;
  signal ptr_deref_936_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_0 : boolean;
  signal ptr_deref_936_store_0_req_1 : boolean;
  signal ptr_deref_936_store_0_ack_1 : boolean;
  signal WPIPE_Block0_start_1000_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1000_inst_req_1 : boolean;
  signal if_stmt_951_branch_req_0 : boolean;
  signal addr_of_1310_final_reg_req_1 : boolean;
  signal if_stmt_951_branch_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_1 : boolean;
  signal if_stmt_951_branch_ack_0 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_ack_1 : boolean;
  signal call_stmt_962_call_req_0 : boolean;
  signal call_stmt_962_call_ack_0 : boolean;
  signal WPIPE_Block1_start_1063_inst_req_1 : boolean;
  signal call_stmt_962_call_req_1 : boolean;
  signal call_stmt_962_call_ack_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_972_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_1 : boolean;
  signal type_cast_1328_inst_ack_1 : boolean;
  signal type_cast_967_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_1 : boolean;
  signal type_cast_967_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_972_inst_req_0 : boolean;
  signal type_cast_967_inst_req_1 : boolean;
  signal type_cast_967_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1000_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_969_inst_req_0 : boolean;
  signal WPIPE_Block0_start_969_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_969_inst_req_1 : boolean;
  signal WPIPE_Block0_start_969_inst_ack_1 : boolean;
  signal array_obj_ref_1309_index_offset_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1390_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1396_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1090_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1090_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1090_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_ack_1 : boolean;
  signal if_stmt_1425_branch_ack_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1093_inst_ack_1 : boolean;
  signal if_stmt_1425_branch_ack_1 : boolean;
  signal type_cast_1318_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1390_inst_ack_0 : boolean;
  signal type_cast_1104_inst_req_0 : boolean;
  signal type_cast_1104_inst_ack_0 : boolean;
  signal type_cast_1104_inst_req_1 : boolean;
  signal type_cast_1104_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1390_inst_req_0 : boolean;
  signal type_cast_1318_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1106_inst_req_0 : boolean;
  signal type_cast_1368_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1106_inst_ack_0 : boolean;
  signal type_cast_1280_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1106_inst_req_1 : boolean;
  signal array_obj_ref_1309_index_offset_req_1 : boolean;
  signal WPIPE_Block2_start_1106_inst_ack_1 : boolean;
  signal type_cast_1111_inst_req_0 : boolean;
  signal type_cast_1368_inst_req_1 : boolean;
  signal type_cast_1111_inst_ack_0 : boolean;
  signal type_cast_1111_inst_req_1 : boolean;
  signal type_cast_1111_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1113_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_req_1 : boolean;
  signal type_cast_1368_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_ack_1 : boolean;
  signal if_stmt_1425_branch_req_0 : boolean;
  signal type_cast_1318_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1116_inst_req_0 : boolean;
  signal type_cast_1368_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1116_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1116_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1116_inst_ack_1 : boolean;
  signal phi_stmt_469_req_0 : boolean;
  signal type_cast_1318_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_0 : boolean;
  signal array_obj_ref_1309_index_offset_ack_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_1 : boolean;
  signal type_cast_1388_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_0 : boolean;
  signal array_obj_ref_1309_index_offset_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_1 : boolean;
  signal type_cast_1388_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1125_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1125_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1125_inst_req_1 : boolean;
  signal type_cast_1358_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1125_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1393_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1128_inst_req_0 : boolean;
  signal type_cast_1358_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1128_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1128_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1128_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1411_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1411_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1393_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_1 : boolean;
  signal type_cast_1358_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_1 : boolean;
  signal type_cast_1388_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_0 : boolean;
  signal type_cast_1358_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1411_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1411_inst_req_0 : boolean;
  signal type_cast_1388_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1399_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1408_inst_ack_1 : boolean;
  signal ptr_deref_1314_load_0_ack_1 : boolean;
  signal ptr_deref_1314_load_0_req_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_1 : boolean;
  signal type_cast_1348_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1408_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1146_inst_req_0 : boolean;
  signal type_cast_1348_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1146_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1146_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1146_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1408_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1408_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_req_1 : boolean;
  signal type_cast_1348_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_ack_1 : boolean;
  signal ptr_deref_1314_load_0_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1399_inst_req_1 : boolean;
  signal type_cast_1160_inst_req_0 : boolean;
  signal type_cast_1348_inst_req_0 : boolean;
  signal type_cast_1160_inst_ack_0 : boolean;
  signal type_cast_1160_inst_req_1 : boolean;
  signal type_cast_1160_inst_ack_1 : boolean;
  signal ptr_deref_1314_load_0_req_0 : boolean;
  signal WPIPE_Block3_start_1162_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1162_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1162_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1162_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1405_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1405_inst_req_1 : boolean;
  signal type_cast_1167_inst_req_0 : boolean;
  signal type_cast_1167_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1399_inst_ack_0 : boolean;
  signal type_cast_1167_inst_req_1 : boolean;
  signal type_cast_1167_inst_ack_1 : boolean;
  signal type_cast_1378_inst_ack_1 : boolean;
  signal type_cast_1378_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1169_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1169_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1169_inst_req_1 : boolean;
  signal type_cast_1338_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1169_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1405_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1405_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1172_inst_req_0 : boolean;
  signal type_cast_1338_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1172_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1172_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1172_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1402_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1402_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_0 : boolean;
  signal type_cast_1338_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_1 : boolean;
  signal type_cast_1338_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1182_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1182_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1182_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1182_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1185_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1185_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1185_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1185_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1188_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1188_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1188_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1188_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1191_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1191_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1191_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1191_inst_ack_1 : boolean;
  signal call_stmt_1195_call_req_0 : boolean;
  signal call_stmt_1195_call_ack_0 : boolean;
  signal call_stmt_1195_call_req_1 : boolean;
  signal call_stmt_1195_call_ack_1 : boolean;
  signal type_cast_1199_inst_req_0 : boolean;
  signal type_cast_1199_inst_ack_0 : boolean;
  signal type_cast_1199_inst_req_1 : boolean;
  signal type_cast_1199_inst_ack_1 : boolean;
  signal type_cast_1208_inst_req_0 : boolean;
  signal type_cast_1208_inst_ack_0 : boolean;
  signal type_cast_1208_inst_req_1 : boolean;
  signal type_cast_1208_inst_ack_1 : boolean;
  signal type_cast_1218_inst_req_0 : boolean;
  signal type_cast_1218_inst_ack_0 : boolean;
  signal type_cast_1218_inst_req_1 : boolean;
  signal type_cast_1218_inst_ack_1 : boolean;
  signal type_cast_1228_inst_req_0 : boolean;
  signal type_cast_1228_inst_ack_0 : boolean;
  signal type_cast_1228_inst_req_1 : boolean;
  signal type_cast_1228_inst_ack_1 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1240_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1240_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1240_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1240_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1243_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1243_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1243_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1243_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1246_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1246_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1246_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1246_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1249_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1249_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1249_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1249_inst_ack_1 : boolean;
  signal if_stmt_1253_branch_req_0 : boolean;
  signal if_stmt_1253_branch_ack_1 : boolean;
  signal if_stmt_1253_branch_ack_0 : boolean;
  signal type_cast_475_inst_req_0 : boolean;
  signal type_cast_475_inst_ack_0 : boolean;
  signal type_cast_475_inst_req_1 : boolean;
  signal type_cast_475_inst_ack_1 : boolean;
  signal phi_stmt_469_req_1 : boolean;
  signal phi_stmt_469_ack_0 : boolean;
  signal phi_stmt_676_req_1 : boolean;
  signal type_cast_679_inst_req_0 : boolean;
  signal type_cast_679_inst_ack_0 : boolean;
  signal type_cast_679_inst_req_1 : boolean;
  signal type_cast_679_inst_ack_1 : boolean;
  signal phi_stmt_676_req_0 : boolean;
  signal phi_stmt_676_ack_0 : boolean;
  signal phi_stmt_920_req_1 : boolean;
  signal type_cast_923_inst_req_0 : boolean;
  signal type_cast_923_inst_ack_0 : boolean;
  signal type_cast_923_inst_req_1 : boolean;
  signal type_cast_923_inst_ack_1 : boolean;
  signal phi_stmt_920_req_0 : boolean;
  signal phi_stmt_920_ack_0 : boolean;
  signal phi_stmt_1297_req_0 : boolean;
  signal type_cast_1303_inst_req_0 : boolean;
  signal type_cast_1303_inst_ack_0 : boolean;
  signal type_cast_1303_inst_req_1 : boolean;
  signal type_cast_1303_inst_ack_1 : boolean;
  signal phi_stmt_1297_req_1 : boolean;
  signal phi_stmt_1297_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(476 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(476);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_32/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/branch_block_stmt_32__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/cr
      -- 
    rr_133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_0); -- 
    cr_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_38_inst_req_1); -- 
    cr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_51_inst_req_1); -- 
    cr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_63_inst_req_1); -- 
    cr_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_76_inst_req_1); -- 
    cr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_88_inst_req_1); -- 
    cr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_101_inst_req_1); -- 
    cr_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_113_inst_req_1); -- 
    cr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_126_inst_req_1); -- 
    cr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_339_inst_req_1); -- 
    cr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_138_inst_req_1); -- 
    cr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_151_inst_req_1); -- 
    cr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_163_inst_req_1); -- 
    cr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_176_inst_req_1); -- 
    cr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_188_inst_req_1); -- 
    cr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_201_inst_req_1); -- 
    cr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_210_inst_req_1); -- 
    cr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_214_inst_req_1); -- 
    cr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_218_inst_req_1); -- 
    cr_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_255_inst_req_1); -- 
    cr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_259_inst_req_1); -- 
    cr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_263_inst_req_1); -- 
    cr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_267_inst_req_1); -- 
    cr_642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_289_inst_req_1); -- 
    cr_670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_302_inst_req_1); -- 
    cr_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_314_inst_req_1); -- 
    cr_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_327_inst_req_1); -- 
    cr_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_352_inst_req_1); -- 
    cr_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_364_inst_req_1); -- 
    cr_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_377_inst_req_1); -- 
    cr_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_389_inst_req_1); -- 
    cr_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_402_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_update_start_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/cr
      -- 
    ra_134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_34_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_sample_start_
      -- 
    ca_139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    rr_147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_38_inst_req_0); -- 
    rr_161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Sample/ra
      -- 
    ra_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_38_Update/ca
      -- 
    ca_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_update_start_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/cr
      -- 
    ra_162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    cr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(5), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_47_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/rr
      -- 
    ca_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    rr_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => type_cast_51_inst_req_0); -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Sample/ra
      -- 
    ra_176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_51_Update/ca
      -- 
    ca_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_update_start_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/cr
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_0, ack => convTranspose_CP_39_elements(9)); -- 
    cr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_59_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/rr
      -- 
    ca_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_1, ack => convTranspose_CP_39_elements(10)); -- 
    rr_203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => type_cast_63_inst_req_0); -- 
    rr_217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Sample/ra
      -- 
    ra_204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_0, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_63_Update/ca
      -- 
    ca_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_1, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_update_start_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/cr
      -- 
    ra_218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_0, ack => convTranspose_CP_39_elements(13)); -- 
    cr_222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(13), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_72_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/rr
      -- 
    ca_223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_1, ack => convTranspose_CP_39_elements(14)); -- 
    rr_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => type_cast_76_inst_req_0); -- 
    rr_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Sample/ra
      -- 
    ra_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => convTranspose_CP_39_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_76_Update/ca
      -- 
    ca_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => convTranspose_CP_39_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_update_start_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/cr
      -- 
    ra_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_84_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/rr
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    rr_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => type_cast_88_inst_req_0); -- 
    rr_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Sample/ra
      -- 
    ra_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_88_Update/ca
      -- 
    ca_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_update_start_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/cr
      -- 
    ra_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_97_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/rr
      -- 
    ca_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_101_inst_req_0); -- 
    rr_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Sample/ra
      -- 
    ra_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_0, ack => convTranspose_CP_39_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_101_Update/ca
      -- 
    ca_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_1, ack => convTranspose_CP_39_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_update_start_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/cr
      -- 
    ra_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_0, ack => convTranspose_CP_39_elements(25)); -- 
    cr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(25), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_109_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/rr
      -- 
    ca_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_1, ack => convTranspose_CP_39_elements(26)); -- 
    rr_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => type_cast_113_inst_req_0); -- 
    rr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Sample/ra
      -- 
    ra_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_0, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_113_Update/ca
      -- 
    ca_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_1, ack => convTranspose_CP_39_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_update_start_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/cr
      -- 
    ra_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_0, ack => convTranspose_CP_39_elements(29)); -- 
    cr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_122_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/rr
      -- 
    ca_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_1, ack => convTranspose_CP_39_elements(30)); -- 
    rr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => type_cast_126_inst_req_0); -- 
    rr_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Sample/ra
      -- 
    ra_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_126_Update/ca
      -- 
    ca_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_update_start_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Sample/ra
      -- 
    ra_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    cr_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(33), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_134_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/rr
      -- 
    ca_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    rr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => type_cast_138_inst_req_0); -- 
    rr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Sample/ra
      -- 
    ra_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_138_Update/ca
      -- 
    ca_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_update_start_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/cr
      -- 
    ra_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_0, ack => convTranspose_CP_39_elements(37)); -- 
    cr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_147_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/rr
      -- 
    ca_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_1, ack => convTranspose_CP_39_elements(38)); -- 
    rr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => type_cast_151_inst_req_0); -- 
    rr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Sample/ra
      -- 
    ra_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_0, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_151_Update/ca
      -- 
    ca_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_1, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_update_start_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/cr
      -- 
    ra_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_0, ack => convTranspose_CP_39_elements(41)); -- 
    cr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(41), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_159_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/rr
      -- 
    ca_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_1, ack => convTranspose_CP_39_elements(42)); -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_0); -- 
    rr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => type_cast_163_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Sample/ra
      -- 
    ra_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_0, ack => convTranspose_CP_39_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_163_Update/ca
      -- 
    ca_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_1, ack => convTranspose_CP_39_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_update_start_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/cr
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    cr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_172_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/rr
      -- 
    ca_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    rr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => type_cast_176_inst_req_0); -- 
    rr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Sample/ra
      -- 
    ra_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_176_Update/ca
      -- 
    ca_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_update_start_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/cr
      -- 
    ra_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_184_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/rr
      -- 
    ca_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_188_inst_req_0); -- 
    rr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Sample/ra
      -- 
    ra_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_0, ack => convTranspose_CP_39_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_188_Update/ca
      -- 
    ca_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_1, ack => convTranspose_CP_39_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_update_start_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/cr
      -- 
    ra_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_0, ack => convTranspose_CP_39_elements(53)); -- 
    cr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(53), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_197_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/rr
      -- 
    ca_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_1, ack => convTranspose_CP_39_elements(54)); -- 
    rr_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => type_cast_201_inst_req_0); -- 
    rr_623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => RPIPE_ConvTranspose_input_pipe_285_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Sample/ra
      -- 
    ra_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_0, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_201_Update/ca
      -- 
    ca_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_1, ack => convTranspose_CP_39_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/rr
      -- 
    rr_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => type_cast_210_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Sample/ra
      -- 
    ra_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_0, ack => convTranspose_CP_39_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_210_Update/ca
      -- 
    ca_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_210_inst_ack_1, ack => convTranspose_CP_39_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/rr
      -- 
    rr_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(60), ack => type_cast_214_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(12) & convTranspose_CP_39_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Sample/ra
      -- 
    ra_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_214_Update/ca
      -- 
    ca_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_214_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/rr
      -- 
    rr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(63), ack => type_cast_218_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(20) & convTranspose_CP_39_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Sample/ra
      -- 
    ra_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_0, ack => convTranspose_CP_39_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_218_Update/ca
      -- 
    ca_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_218_inst_ack_1, ack => convTranspose_CP_39_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/rr
      -- 
    rr_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => type_cast_255_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(28) & convTranspose_CP_39_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Sample/ra
      -- 
    ra_568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_0, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_255_Update/ca
      -- 
    ca_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_1, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/rr
      -- 
    rr_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(69), ack => type_cast_259_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(40) & convTranspose_CP_39_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Sample/ra
      -- 
    ra_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_259_inst_ack_0, ack => convTranspose_CP_39_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_259_Update/ca
      -- 
    ca_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_259_inst_ack_1, ack => convTranspose_CP_39_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	44 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/rr
      -- 
    rr_595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(72), ack => type_cast_263_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(44) & convTranspose_CP_39_elements(48);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Sample/ra
      -- 
    ra_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_263_Update/ca
      -- 
    ca_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: 	56 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/rr
      -- 
    rr_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(75), ack => type_cast_267_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(52) & convTranspose_CP_39_elements(56);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Sample/ra
      -- 
    ra_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_0, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_267_Update/ca
      -- 
    ca_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_1, ack => convTranspose_CP_39_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_update_start_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/cr
      -- 
    ra_624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_285_inst_ack_0, ack => convTranspose_CP_39_elements(78)); -- 
    cr_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_285_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_285_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/rr
      -- 
    ca_629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_285_inst_ack_1, ack => convTranspose_CP_39_elements(79)); -- 
    rr_637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => type_cast_289_inst_req_0); -- 
    rr_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(79), ack => RPIPE_ConvTranspose_input_pipe_298_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Sample/ra
      -- 
    ra_638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_289_inst_ack_0, ack => convTranspose_CP_39_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_289_Update/ca
      -- 
    ca_643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_289_inst_ack_1, ack => convTranspose_CP_39_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_update_start_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/cr
      -- 
    ra_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_298_inst_ack_0, ack => convTranspose_CP_39_elements(82)); -- 
    cr_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => RPIPE_ConvTranspose_input_pipe_298_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_298_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/rr
      -- 
    ca_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_298_inst_ack_1, ack => convTranspose_CP_39_elements(83)); -- 
    rr_665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => type_cast_302_inst_req_0); -- 
    rr_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(83), ack => RPIPE_ConvTranspose_input_pipe_310_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Sample/ra
      -- 
    ra_666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_0, ack => convTranspose_CP_39_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_302_Update/ca
      -- 
    ca_671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_302_inst_ack_1, ack => convTranspose_CP_39_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_update_start_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/cr
      -- 
    ra_680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_310_inst_ack_0, ack => convTranspose_CP_39_elements(86)); -- 
    cr_684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => RPIPE_ConvTranspose_input_pipe_310_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_310_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/rr
      -- 
    ca_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_310_inst_ack_1, ack => convTranspose_CP_39_elements(87)); -- 
    rr_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => type_cast_314_inst_req_0); -- 
    rr_707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(87), ack => RPIPE_ConvTranspose_input_pipe_323_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Sample/ra
      -- 
    ra_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_314_inst_ack_0, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_314_Update/ca
      -- 
    ca_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_314_inst_ack_1, ack => convTranspose_CP_39_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_update_start_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/cr
      -- 
    ra_708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_323_inst_ack_0, ack => convTranspose_CP_39_elements(90)); -- 
    cr_712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => RPIPE_ConvTranspose_input_pipe_323_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_323_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/rr
      -- 
    ca_713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_323_inst_ack_1, ack => convTranspose_CP_39_elements(91)); -- 
    rr_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => type_cast_327_inst_req_0); -- 
    rr_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(91), ack => RPIPE_ConvTranspose_input_pipe_335_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Sample/ra
      -- 
    ra_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_327_inst_ack_0, ack => convTranspose_CP_39_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_327_Update/ca
      -- 
    ca_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_327_inst_ack_1, ack => convTranspose_CP_39_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_update_start_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/cr
      -- 
    ra_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_335_inst_ack_0, ack => convTranspose_CP_39_elements(94)); -- 
    cr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(94), ack => RPIPE_ConvTranspose_input_pipe_335_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_335_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/$entry
      -- 
    ca_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_335_inst_ack_1, ack => convTranspose_CP_39_elements(95)); -- 
    rr_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => type_cast_339_inst_req_0); -- 
    rr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(95), ack => RPIPE_ConvTranspose_input_pipe_348_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Sample/$exit
      -- 
    ra_750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_339_inst_ack_0, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_339_update_completed_
      -- 
    ca_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_339_inst_ack_1, ack => convTranspose_CP_39_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_update_start_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/cr
      -- 
    ra_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_348_inst_ack_0, ack => convTranspose_CP_39_elements(98)); -- 
    cr_768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => RPIPE_ConvTranspose_input_pipe_348_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_348_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/rr
      -- 
    ca_769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_348_inst_ack_1, ack => convTranspose_CP_39_elements(99)); -- 
    rr_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => type_cast_352_inst_req_0); -- 
    rr_791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(99), ack => RPIPE_ConvTranspose_input_pipe_360_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Sample/ra
      -- 
    ra_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_352_inst_ack_0, ack => convTranspose_CP_39_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_352_Update/ca
      -- 
    ca_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_352_inst_ack_1, ack => convTranspose_CP_39_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_update_start_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/cr
      -- 
    ra_792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_360_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    cr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(102), ack => RPIPE_ConvTranspose_input_pipe_360_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_360_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/rr
      -- 
    ca_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_360_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    rr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => type_cast_364_inst_req_0); -- 
    rr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(103), ack => RPIPE_ConvTranspose_input_pipe_373_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Sample/ra
      -- 
    ra_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_364_inst_ack_0, ack => convTranspose_CP_39_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_364_Update/ca
      -- 
    ca_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_364_inst_ack_1, ack => convTranspose_CP_39_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_update_start_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/cr
      -- 
    ra_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_373_inst_ack_0, ack => convTranspose_CP_39_elements(106)); -- 
    cr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(106), ack => RPIPE_ConvTranspose_input_pipe_373_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_373_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/rr
      -- 
    ca_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_373_inst_ack_1, ack => convTranspose_CP_39_elements(107)); -- 
    rr_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => type_cast_377_inst_req_0); -- 
    rr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(107), ack => RPIPE_ConvTranspose_input_pipe_385_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Sample/ra
      -- 
    ra_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_377_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_377_Update/ca
      -- 
    ca_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_377_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_update_start_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/cr
      -- 
    ra_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_385_inst_ack_0, ack => convTranspose_CP_39_elements(110)); -- 
    cr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(110), ack => RPIPE_ConvTranspose_input_pipe_385_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_385_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/rr
      -- 
    ca_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_385_inst_ack_1, ack => convTranspose_CP_39_elements(111)); -- 
    rr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => type_cast_389_inst_req_0); -- 
    rr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(111), ack => RPIPE_ConvTranspose_input_pipe_398_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Sample/ra
      -- 
    ra_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_389_inst_ack_0, ack => convTranspose_CP_39_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_389_Update/ca
      -- 
    ca_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_389_inst_ack_1, ack => convTranspose_CP_39_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_update_start_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/cr
      -- 
    ra_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_398_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    cr_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(114), ack => RPIPE_ConvTranspose_input_pipe_398_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/RPIPE_ConvTranspose_input_pipe_398_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/rr
      -- 
    ca_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_398_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    rr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(115), ack => type_cast_402_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Sample/ra
      -- 
    ra_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_402_inst_ack_0, ack => convTranspose_CP_39_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/type_cast_402_Update/ca
      -- 
    ca_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_402_inst_ack_1, ack => convTranspose_CP_39_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415__exit__
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416__entry__
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_415/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_32/R_cmp505_417_place
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/if_stmt_416_else_link/$entry
      -- 
    branch_req_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(118), ack => if_stmt_416_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(65) & convTranspose_CP_39_elements(68) & convTranspose_CP_39_elements(62) & convTranspose_CP_39_elements(59) & convTranspose_CP_39_elements(71) & convTranspose_CP_39_elements(74) & convTranspose_CP_39_elements(77) & convTranspose_CP_39_elements(81) & convTranspose_CP_39_elements(85) & convTranspose_CP_39_elements(89) & convTranspose_CP_39_elements(93) & convTranspose_CP_39_elements(97) & convTranspose_CP_39_elements(101) & convTranspose_CP_39_elements(105) & convTranspose_CP_39_elements(109) & convTranspose_CP_39_elements(113) & convTranspose_CP_39_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437__exit__
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466__entry__
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_416_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_416_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph507
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_update_start_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiAck/dummy
      -- CP-element group 119: 	 branch_block_stmt_32/merge_stmt_437_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph507_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/entry_bbx_xnph507_PhiReq/$entry
      -- 
    if_choice_transition_908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_416_branch_ack_1, ack => convTranspose_CP_39_elements(119)); -- 
    rr_947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_452_inst_req_0); -- 
    cr_952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(119), ack => type_cast_452_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	449 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_416_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_416_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- 
    else_choice_transition_912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_416_branch_ack_0, ack => convTranspose_CP_39_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	449 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638__exit__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673__entry__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_update_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_431_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_431_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph503
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph503_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph503_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_638_PhiAck/dummy
      -- 
    if_choice_transition_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_431_branch_ack_1, ack => convTranspose_CP_39_elements(121)); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_659_inst_req_1); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_659_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	449 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	462 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_431_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_431_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_431_branch_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Sample/ra
      -- 
    ra_948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_0, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	450 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466__exit__
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_443_to_assign_stmt_466/type_cast_452_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody_PhiReq/phi_stmt_469/$entry
      -- CP-element group 124: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody_PhiReq/$entry
      -- 
    ca_953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_452_inst_ack_1, ack => convTranspose_CP_39_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	455 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/ack
      -- 
    ack_982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_481_index_offset_ack_0, ack => convTranspose_CP_39_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	455 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/req
      -- 
    ack_987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_481_index_offset_ack_1, ack => convTranspose_CP_39_elements(126)); -- 
    req_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(126), ack => addr_of_482_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_request/ack
      -- 
    ack_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_482_final_reg_ack_0, ack => convTranspose_CP_39_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	455 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/ack
      -- 
    ack_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_482_final_reg_ack_1, ack => convTranspose_CP_39_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	455 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_update_start_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/cr
      -- 
    ra_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_485_inst_ack_0, ack => convTranspose_CP_39_elements(129)); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => RPIPE_ConvTranspose_input_pipe_485_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/rr
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_485_inst_ack_1, ack => convTranspose_CP_39_elements(130)); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => type_cast_489_inst_req_0); -- 
    rr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(130), ack => RPIPE_ConvTranspose_input_pipe_498_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Sample/ra
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_489_inst_ack_0, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	455 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/ca
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_489_inst_ack_1, ack => convTranspose_CP_39_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_update_start_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/cr
      -- 
    ra_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_498_inst_ack_0, ack => convTranspose_CP_39_elements(133)); -- 
    cr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => RPIPE_ConvTranspose_input_pipe_498_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_498_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/rr
      -- 
    ca_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_498_inst_ack_1, ack => convTranspose_CP_39_elements(134)); -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => type_cast_502_inst_req_0); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(134), ack => RPIPE_ConvTranspose_input_pipe_516_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Sample/ra
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_502_inst_ack_0, ack => convTranspose_CP_39_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	455 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/ca
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_502_inst_ack_1, ack => convTranspose_CP_39_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_update_start_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/cr
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_516_inst_ack_0, ack => convTranspose_CP_39_elements(137)); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => RPIPE_ConvTranspose_input_pipe_516_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_516_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_sample_start_
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_516_inst_ack_1, ack => convTranspose_CP_39_elements(138)); -- 
    rr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => type_cast_520_inst_req_0); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(138), ack => RPIPE_ConvTranspose_input_pipe_534_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Sample/ra
      -- 
    ra_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_0, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	455 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/ca
      -- 
    ca_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_1, ack => convTranspose_CP_39_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_update_start_
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_534_inst_ack_0, ack => convTranspose_CP_39_elements(141)); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => RPIPE_ConvTranspose_input_pipe_534_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_534_update_completed_
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_534_inst_ack_1, ack => convTranspose_CP_39_elements(142)); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => type_cast_538_inst_req_0); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(142), ack => RPIPE_ConvTranspose_input_pipe_552_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_sample_completed_
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_0, ack => convTranspose_CP_39_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	455 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/$exit
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_1, ack => convTranspose_CP_39_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_update_start_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Sample/$exit
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_552_inst_ack_0, ack => convTranspose_CP_39_elements(145)); -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => RPIPE_ConvTranspose_input_pipe_552_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_552_Update/$exit
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_552_inst_ack_1, ack => convTranspose_CP_39_elements(146)); -- 
    rr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => type_cast_556_inst_req_0); -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(146), ack => RPIPE_ConvTranspose_input_pipe_570_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_sample_completed_
      -- 
    ra_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_556_inst_ack_0, ack => convTranspose_CP_39_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	455 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_update_completed_
      -- 
    ca_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_556_inst_ack_1, ack => convTranspose_CP_39_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_update_start_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_sample_completed_
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_570_inst_ack_0, ack => convTranspose_CP_39_elements(149)); -- 
    cr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => RPIPE_ConvTranspose_input_pipe_570_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_570_update_completed_
      -- 
    ca_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_570_inst_ack_1, ack => convTranspose_CP_39_elements(150)); -- 
    rr_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => type_cast_574_inst_req_0); -- 
    rr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(150), ack => RPIPE_ConvTranspose_input_pipe_588_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_sample_completed_
      -- 
    ra_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_0, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	455 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_update_completed_
      -- 
    ca_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_1, ack => convTranspose_CP_39_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_update_start_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_sample_completed_
      -- 
    ra_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_588_inst_ack_0, ack => convTranspose_CP_39_elements(153)); -- 
    cr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => RPIPE_ConvTranspose_input_pipe_588_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_588_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_sample_start_
      -- 
    ca_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_588_inst_ack_1, ack => convTranspose_CP_39_elements(154)); -- 
    rr_1192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => type_cast_592_inst_req_0); -- 
    rr_1206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(154), ack => RPIPE_ConvTranspose_input_pipe_606_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_sample_completed_
      -- 
    ra_1193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_0, ack => convTranspose_CP_39_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	455 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/ca
      -- 
    ca_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_1, ack => convTranspose_CP_39_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_update_start_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_sample_completed_
      -- 
    ra_1207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_606_inst_ack_0, ack => convTranspose_CP_39_elements(157)); -- 
    cr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => RPIPE_ConvTranspose_input_pipe_606_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_606_update_completed_
      -- 
    ca_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_606_inst_ack_1, ack => convTranspose_CP_39_elements(158)); -- 
    rr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(158), ack => type_cast_610_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_sample_completed_
      -- 
    ra_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_0, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	455 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_update_completed_
      -- 
    ca_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_610_inst_ack_1, ack => convTranspose_CP_39_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/ptr_deref_618_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/$entry
      -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => ptr_deref_618_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(128) & convTranspose_CP_39_elements(132) & convTranspose_CP_39_elements(136) & convTranspose_CP_39_elements(140) & convTranspose_CP_39_elements(144) & convTranspose_CP_39_elements(148) & convTranspose_CP_39_elements(152) & convTranspose_CP_39_elements(156) & convTranspose_CP_39_elements(160);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Sample/$exit
      -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_618_store_0_ack_0, ack => convTranspose_CP_39_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	455 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_update_completed_
      -- 
    ca_1276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_618_store_0_ack_1, ack => convTranspose_CP_39_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631__exit__
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632__entry__
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/R_exitcond3_633_place
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/if_stmt_632_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/$exit
      -- 
    branch_req_1284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => if_stmt_632_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(163) & convTranspose_CP_39_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	449 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_632_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422__exit__
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_632_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/merge_stmt_422_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- 
    if_choice_transition_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_632_branch_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	451 
    -- CP-element group 166: 	452 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_632_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_632_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_632_branch_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    rr_3394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_475_inst_req_0); -- 
    cr_3399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(166), ack => type_cast_475_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_sample_completed_
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_0, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	456 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673__exit__
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph503_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/type_cast_659_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_644_to_assign_stmt_673/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph503_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph503_forx_xbody196_PhiReq/phi_stmt_676/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/bbx_xnph503_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$entry
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_1, ack => convTranspose_CP_39_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	461 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_sample_complete
      -- 
    ack_1341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_688_index_offset_ack_0, ack => convTranspose_CP_39_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	461 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/req
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_base_plus_offset/sum_rename_ack
      -- 
    ack_1346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_688_index_offset_ack_1, ack => convTranspose_CP_39_elements(170)); -- 
    req_1355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(170), ack => addr_of_689_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/ack
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_request/$exit
      -- 
    ack_1356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_689_final_reg_ack_0, ack => convTranspose_CP_39_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	461 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_word_addrgen/root_register_ack
      -- 
    ack_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_689_final_reg_ack_1, ack => convTranspose_CP_39_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	461 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_update_start_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/$exit
      -- 
    ra_1370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_692_inst_ack_0, ack => convTranspose_CP_39_elements(173)); -- 
    cr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => RPIPE_ConvTranspose_input_pipe_692_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_sample_start_
      -- 
    ca_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_692_inst_ack_1, ack => convTranspose_CP_39_elements(174)); -- 
    rr_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => type_cast_696_inst_req_0); -- 
    rr_1397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(174), ack => RPIPE_ConvTranspose_input_pipe_705_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_sample_completed_
      -- 
    ra_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_696_inst_ack_0, ack => convTranspose_CP_39_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	461 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_update_completed_
      -- 
    ca_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_696_inst_ack_1, ack => convTranspose_CP_39_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_update_start_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_sample_completed_
      -- 
    ra_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_705_inst_ack_0, ack => convTranspose_CP_39_elements(177)); -- 
    cr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => RPIPE_ConvTranspose_input_pipe_705_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_705_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_sample_start_
      -- 
    ca_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_705_inst_ack_1, ack => convTranspose_CP_39_elements(178)); -- 
    rr_1411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => type_cast_709_inst_req_0); -- 
    rr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(178), ack => RPIPE_ConvTranspose_input_pipe_723_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Sample/$exit
      -- 
    ra_1412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_0, ack => convTranspose_CP_39_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	461 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/$exit
      -- 
    ca_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_1, ack => convTranspose_CP_39_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_update_start_
      -- 
    ra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_723_inst_ack_0, ack => convTranspose_CP_39_elements(181)); -- 
    cr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => RPIPE_ConvTranspose_input_pipe_723_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_723_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_sample_start_
      -- 
    ca_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_723_inst_ack_1, ack => convTranspose_CP_39_elements(182)); -- 
    rr_1439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => type_cast_727_inst_req_0); -- 
    rr_1453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => RPIPE_ConvTranspose_input_pipe_741_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_sample_completed_
      -- 
    ra_1440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_0, ack => convTranspose_CP_39_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	461 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_update_completed_
      -- 
    ca_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_1, ack => convTranspose_CP_39_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/cr
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_update_start_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Sample/ra
      -- 
    ra_1454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_741_inst_ack_0, ack => convTranspose_CP_39_elements(185)); -- 
    cr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(185), ack => RPIPE_ConvTranspose_input_pipe_741_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	189 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_741_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/rr
      -- 
    ca_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_741_inst_ack_1, ack => convTranspose_CP_39_elements(186)); -- 
    rr_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => RPIPE_ConvTranspose_input_pipe_759_inst_req_0); -- 
    rr_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(186), ack => type_cast_745_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Sample/ra
      -- 
    ra_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_745_inst_ack_0, ack => convTranspose_CP_39_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	461 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/ca
      -- 
    ca_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_745_inst_ack_1, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_update_start_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/cr
      -- 
    ra_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_759_inst_ack_0, ack => convTranspose_CP_39_elements(189)); -- 
    cr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => RPIPE_ConvTranspose_input_pipe_759_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	193 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_759_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/rr
      -- 
    ca_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_759_inst_ack_1, ack => convTranspose_CP_39_elements(190)); -- 
    rr_1495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_763_inst_req_0); -- 
    rr_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => RPIPE_ConvTranspose_input_pipe_777_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Sample/ra
      -- 
    ra_1496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_0, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	461 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/ca
      -- 
    ca_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_763_inst_ack_1, ack => convTranspose_CP_39_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_update_start_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/cr
      -- 
    ra_1510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_777_inst_ack_0, ack => convTranspose_CP_39_elements(193)); -- 
    cr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(193), ack => RPIPE_ConvTranspose_input_pipe_777_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_777_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/rr
      -- 
    ca_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_777_inst_ack_1, ack => convTranspose_CP_39_elements(194)); -- 
    rr_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => type_cast_781_inst_req_0); -- 
    rr_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => RPIPE_ConvTranspose_input_pipe_795_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Sample/ra
      -- 
    ra_1524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_0, ack => convTranspose_CP_39_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	461 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/ca
      -- 
    ca_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_1, ack => convTranspose_CP_39_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_update_start_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/cr
      -- 
    ra_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_795_inst_ack_0, ack => convTranspose_CP_39_elements(197)); -- 
    cr_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(197), ack => RPIPE_ConvTranspose_input_pipe_795_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_795_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/rr
      -- 
    ca_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_795_inst_ack_1, ack => convTranspose_CP_39_elements(198)); -- 
    rr_1551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => type_cast_799_inst_req_0); -- 
    rr_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(198), ack => RPIPE_ConvTranspose_input_pipe_813_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Sample/ra
      -- 
    ra_1552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_0, ack => convTranspose_CP_39_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	461 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/ca
      -- 
    ca_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_1, ack => convTranspose_CP_39_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_update_start_
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/cr
      -- 
    ra_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_813_inst_ack_0, ack => convTranspose_CP_39_elements(201)); -- 
    cr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => RPIPE_ConvTranspose_input_pipe_813_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_813_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/rr
      -- 
    ca_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_813_inst_ack_1, ack => convTranspose_CP_39_elements(202)); -- 
    rr_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => type_cast_817_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Sample/ra
      -- 
    ra_1580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_0, ack => convTranspose_CP_39_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	461 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/ca
      -- 
    ca_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_1, ack => convTranspose_CP_39_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/ptr_deref_825_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/rr
      -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(205), ack => ptr_deref_825_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(196) & convTranspose_CP_39_elements(200) & convTranspose_CP_39_elements(204) & convTranspose_CP_39_elements(192) & convTranspose_CP_39_elements(172) & convTranspose_CP_39_elements(176) & convTranspose_CP_39_elements(180) & convTranspose_CP_39_elements(184) & convTranspose_CP_39_elements(188);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Sample/word_access_start/word_0/ra
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_825_store_0_ack_0, ack => convTranspose_CP_39_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	461 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/ca
      -- 
    ca_1635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_825_store_0_ack_1, ack => convTranspose_CP_39_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	169 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838__exit__
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839__entry__
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_32/R_exitcond2_840_place
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/if_stmt_839_else_link/$entry
      -- 
    branch_req_1643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => if_stmt_839_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(207) & convTranspose_CP_39_elements(169);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	462 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845__exit__
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_839_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_839_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/merge_stmt_845_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_839_branch_ack_1, ack => convTranspose_CP_39_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	457 
    -- CP-element group 210: 	458 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_839_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_839_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_839_branch_ack_0, ack => convTranspose_CP_39_elements(210)); -- 
    rr_3448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_679_inst_req_0); -- 
    cr_3453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => type_cast_679_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	462 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/ra
      -- 
    ra_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	462 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/ca
      -- 
    ca_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	462 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/ra
      -- 
    ra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	462 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/ca
      -- 
    ca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	462 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/ra
      -- 
    ra_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_858_inst_ack_0, ack => convTranspose_CP_39_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	462 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/ca
      -- 
    ca_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_858_inst_ack_1, ack => convTranspose_CP_39_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875__exit__
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876__entry__
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_32/R_cmp264497_877_place
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_876_else_link/$entry
      -- 
    branch_req_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(217), ack => if_stmt_876_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(212) & convTranspose_CP_39_elements(214) & convTranspose_CP_39_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882__exit__
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917__entry__
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_876_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_876_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph499
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_update_start_
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph499_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend250_bbx_xnph499_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_882_PhiAck/dummy
      -- 
    if_choice_transition_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_876_branch_ack_1, ack => convTranspose_CP_39_elements(218)); -- 
    rr_1729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_903_inst_req_0); -- 
    cr_1734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => type_cast_903_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	469 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_876_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_876_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_876_branch_ack_0, ack => convTranspose_CP_39_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Sample/ra
      -- 
    ra_1730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_0, ack => convTranspose_CP_39_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	463 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917__exit__
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph499_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_888_to_assign_stmt_917/type_cast_903_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph499_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph499_forx_xbody266_PhiReq/phi_stmt_920/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/bbx_xnph499_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$entry
      -- 
    ca_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_1, ack => convTranspose_CP_39_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	468 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/ack
      -- 
    ack_1764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_offset_ack_0, ack => convTranspose_CP_39_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	468 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/req
      -- 
    ack_1769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_932_index_offset_ack_1, ack => convTranspose_CP_39_elements(223)); -- 
    req_1778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => addr_of_933_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_request/ack
      -- 
    ack_1779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_933_final_reg_ack_0, ack => convTranspose_CP_39_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	468 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/ptr_deref_936_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/rr
      -- 
    ack_1784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_933_final_reg_ack_1, ack => convTranspose_CP_39_elements(225)); -- 
    rr_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(225), ack => ptr_deref_936_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Sample/word_access_start/word_0/ra
      -- 
    ra_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_936_store_0_ack_0, ack => convTranspose_CP_39_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	468 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/ca
      -- 
    ca_1834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_936_store_0_ack_1, ack => convTranspose_CP_39_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950__exit__
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951__entry__
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_32/R_exitcond_952_place
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/if_stmt_951_else_link/$entry
      -- 
    branch_req_1842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => if_stmt_951_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(222) & convTranspose_CP_39_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	469 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957__exit__
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_951_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_951_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/merge_stmt_957_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_951_branch_ack_1, ack => convTranspose_CP_39_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	464 
    -- CP-element group 230: 	465 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_32/if_stmt_951_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/if_stmt_951_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_951_branch_ack_0, ack => convTranspose_CP_39_elements(230)); -- 
    rr_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_923_inst_req_0); -- 
    cr_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => type_cast_923_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	469 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Sample/cra
      -- 
    cra_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_962_call_ack_0, ack => convTranspose_CP_39_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	469 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Sample/rr
      -- 
    cca_1870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_962_call_ack_1, ack => convTranspose_CP_39_elements(232)); -- 
    rr_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(232), ack => type_cast_967_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Sample/ra
      -- 
    ra_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_0, ack => convTranspose_CP_39_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	469 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	373 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Update/ca
      -- 
    ca_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_1, ack => convTranspose_CP_39_elements(234)); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	469 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_update_start_
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Update/req
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_969_inst_ack_0, ack => convTranspose_CP_39_elements(235)); -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => WPIPE_Block0_start_969_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Sample/req
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Sample/$entry
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_969_inst_ack_1, ack => convTranspose_CP_39_elements(236)); -- 
    req_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_Block0_start_972_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Update/req
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_update_start_
      -- 
    ack_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_972_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_Block0_start_972_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Sample/req
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_972_update_completed_
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_972_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(238), ack => WPIPE_Block0_start_975_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_update_start_
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Update/req
      -- 
    ack_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    req_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(239), ack => WPIPE_Block0_start_975_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_975_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Sample/req
      -- 
    ack_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    req_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(240), ack => WPIPE_Block0_start_978_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Update/req
      -- 
    ack_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => WPIPE_Block0_start_978_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Sample/req
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_978_Update/ack
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    req_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => WPIPE_Block0_start_981_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Update/req
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_update_start_
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_sample_completed_
      -- 
    ack_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_0, ack => convTranspose_CP_39_elements(243)); -- 
    req_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_Block0_start_981_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_981_update_completed_
      -- 
    ack_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_1, ack => convTranspose_CP_39_elements(244)); -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_Block0_start_984_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Update/req
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_update_start_
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_sample_completed_
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_0, ack => convTranspose_CP_39_elements(245)); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(245), ack => WPIPE_Block0_start_984_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_984_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Sample/$entry
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_1, ack => convTranspose_CP_39_elements(246)); -- 
    req_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(246), ack => WPIPE_Block0_start_987_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Update/req
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_update_start_
      -- 
    ack_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_0, ack => convTranspose_CP_39_elements(247)); -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(247), ack => WPIPE_Block0_start_987_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Sample/req
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_987_update_completed_
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_1, ack => convTranspose_CP_39_elements(248)); -- 
    req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => WPIPE_Block0_start_990_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Update/req
      -- 
    ack_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_0, ack => convTranspose_CP_39_elements(249)); -- 
    req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => WPIPE_Block0_start_990_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_990_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Sample/req
      -- 
    ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_1, ack => convTranspose_CP_39_elements(250)); -- 
    req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_Block0_start_993_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_update_start_
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Update/req
      -- 
    ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_Block0_start_993_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_993_Update/ack
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    req_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(252), ack => WPIPE_Block0_start_996_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Update/req
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_update_start_
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_sample_completed_
      -- 
    ack_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_996_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    req_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(253), ack => WPIPE_Block0_start_996_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Sample/req
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_996_update_completed_
      -- 
    ack_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_996_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    req_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(254), ack => WPIPE_Block0_start_1000_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Update/req
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Sample/ack
      -- 
    ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1000_inst_ack_0, ack => convTranspose_CP_39_elements(255)); -- 
    req_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => WPIPE_Block0_start_1000_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1000_Update/$exit
      -- 
    ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1000_inst_ack_1, ack => convTranspose_CP_39_elements(256)); -- 
    req_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(256), ack => WPIPE_Block0_start_1004_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Update/req
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_update_start_
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_sample_completed_
      -- 
    ack_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1004_inst_ack_0, ack => convTranspose_CP_39_elements(257)); -- 
    req_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(257), ack => WPIPE_Block0_start_1004_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Sample/req
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1004_update_completed_
      -- 
    ack_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1004_inst_ack_1, ack => convTranspose_CP_39_elements(258)); -- 
    req_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(258), ack => WPIPE_Block0_start_1007_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Update/req
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_sample_completed_
      -- 
    ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1007_inst_ack_0, ack => convTranspose_CP_39_elements(259)); -- 
    req_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(259), ack => WPIPE_Block0_start_1007_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1007_update_completed_
      -- 
    ack_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1007_inst_ack_1, ack => convTranspose_CP_39_elements(260)); -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => WPIPE_Block0_start_1010_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Update/req
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_update_start_
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_sample_completed_
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1010_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    req_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(261), ack => WPIPE_Block0_start_1010_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	373 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_1010_update_completed_
      -- 
    ack_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1010_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	469 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_update_start_
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Update/req
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_sample_completed_
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1013_inst_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(263), ack => WPIPE_Block1_start_1013_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Sample/req
      -- 
    ack_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1013_inst_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    req_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => WPIPE_Block1_start_1016_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Update/req
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_update_start_
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Update/$entry
      -- 
    ack_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1016_inst_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    req_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(265), ack => WPIPE_Block1_start_1016_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1016_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Sample/req
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_sample_start_
      -- 
    ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1016_inst_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    req_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(266), ack => WPIPE_Block1_start_1019_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Update/req
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_update_start_
      -- 
    ack_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(267), ack => WPIPE_Block1_start_1019_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1019_update_completed_
      -- 
    ack_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    req_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => WPIPE_Block1_start_1022_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Update/req
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_update_start_
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_sample_completed_
      -- 
    ack_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(269), ack => WPIPE_Block1_start_1022_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1022_update_completed_
      -- 
    ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    req_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(270), ack => WPIPE_Block1_start_1025_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_update_start_
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Update/req
      -- 
    ack_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(271), ack => WPIPE_Block1_start_1025_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1025_Update/$exit
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    req_2158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(272), ack => WPIPE_Block1_start_1028_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Update/req
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_update_start_
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_sample_completed_
      -- 
    ack_2159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    req_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(273), ack => WPIPE_Block1_start_1028_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1028_update_completed_
      -- 
    ack_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    req_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => WPIPE_Block1_start_1031_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Update/req
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_sample_completed_
      -- 
    ack_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_0, ack => convTranspose_CP_39_elements(275)); -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(275), ack => WPIPE_Block1_start_1031_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1031_update_completed_
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_1, ack => convTranspose_CP_39_elements(276)); -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(276), ack => WPIPE_Block1_start_1034_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Update/req
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_update_start_
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_sample_completed_
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1034_inst_ack_0, ack => convTranspose_CP_39_elements(277)); -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(277), ack => WPIPE_Block1_start_1034_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1034_update_completed_
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1034_inst_ack_1, ack => convTranspose_CP_39_elements(278)); -- 
    req_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(278), ack => WPIPE_Block1_start_1037_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Update/req
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_update_start_
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_sample_completed_
      -- 
    ack_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_0, ack => convTranspose_CP_39_elements(279)); -- 
    req_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(279), ack => WPIPE_Block1_start_1037_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1037_update_completed_
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_1, ack => convTranspose_CP_39_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	469 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Sample/ra
      -- 
    ra_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1048_inst_ack_0, ack => convTranspose_CP_39_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	469 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Update/ca
      -- 
    ca_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1048_inst_ack_1, ack => convTranspose_CP_39_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	280 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Sample/req
      -- 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(283), ack => WPIPE_Block1_start_1050_inst_req_0); -- 
    convTranspose_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(280) & convTranspose_CP_39_elements(282);
      gj_convTranspose_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_update_start_
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Update/req
      -- 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1050_inst_ack_0, ack => convTranspose_CP_39_elements(284)); -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(284), ack => WPIPE_Block1_start_1050_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	288 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1050_Update/ack
      -- 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1050_inst_ack_1, ack => convTranspose_CP_39_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	469 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Sample/ra
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_sample_completed_
      -- 
    ra_2243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_0, ack => convTranspose_CP_39_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	469 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_update_completed_
      -- 
    ca_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_1, ack => convTranspose_CP_39_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_sample_start_
      -- 
    req_2256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => WPIPE_Block1_start_1057_inst_req_0); -- 
    convTranspose_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(285) & convTranspose_CP_39_elements(287);
      gj_convTranspose_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Update/req
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_sample_completed_
      -- 
    ack_2257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1057_inst_ack_0, ack => convTranspose_CP_39_elements(289)); -- 
    req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(289), ack => WPIPE_Block1_start_1057_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1057_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_sample_start_
      -- 
    ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1057_inst_ack_1, ack => convTranspose_CP_39_elements(290)); -- 
    req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(290), ack => WPIPE_Block1_start_1060_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Update/req
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_update_start_
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_sample_completed_
      -- 
    ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1060_inst_ack_0, ack => convTranspose_CP_39_elements(291)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(291), ack => WPIPE_Block1_start_1060_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1060_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Sample/$entry
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1060_inst_ack_1, ack => convTranspose_CP_39_elements(292)); -- 
    req_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(292), ack => WPIPE_Block1_start_1063_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Update/req
      -- 
    ack_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1063_inst_ack_0, ack => convTranspose_CP_39_elements(293)); -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(293), ack => WPIPE_Block1_start_1063_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1063_Update/$exit
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1063_inst_ack_1, ack => convTranspose_CP_39_elements(294)); -- 
    req_2298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => WPIPE_Block1_start_1066_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Update/req
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_sample_completed_
      -- 
    ack_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1066_inst_ack_0, ack => convTranspose_CP_39_elements(295)); -- 
    req_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(295), ack => WPIPE_Block1_start_1066_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	373 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1066_update_completed_
      -- 
    ack_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1066_inst_ack_1, ack => convTranspose_CP_39_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	469 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_update_start_
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Update/req
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Sample/$exit
      -- 
    ack_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1069_inst_ack_0, ack => convTranspose_CP_39_elements(297)); -- 
    req_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(297), ack => WPIPE_Block2_start_1069_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Sample/$entry
      -- 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1069_inst_ack_1, ack => convTranspose_CP_39_elements(298)); -- 
    req_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(298), ack => WPIPE_Block2_start_1072_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Update/req
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_update_start_
      -- 
    ack_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1072_inst_ack_0, ack => convTranspose_CP_39_elements(299)); -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(299), ack => WPIPE_Block2_start_1072_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1072_update_completed_
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1072_inst_ack_1, ack => convTranspose_CP_39_elements(300)); -- 
    req_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(300), ack => WPIPE_Block2_start_1075_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Update/req
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Sample/$exit
      -- 
    ack_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_0, ack => convTranspose_CP_39_elements(301)); -- 
    req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(301), ack => WPIPE_Block2_start_1075_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1075_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_sample_start_
      -- 
    ack_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_1, ack => convTranspose_CP_39_elements(302)); -- 
    req_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => WPIPE_Block2_start_1078_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Update/req
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_update_start_
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_sample_completed_
      -- 
    ack_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_0, ack => convTranspose_CP_39_elements(303)); -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(303), ack => WPIPE_Block2_start_1078_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1078_update_completed_
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_1, ack => convTranspose_CP_39_elements(304)); -- 
    req_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(304), ack => WPIPE_Block2_start_1081_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Update/req
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_update_start_
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Sample/ack
      -- 
    ack_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_0, ack => convTranspose_CP_39_elements(305)); -- 
    req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(305), ack => WPIPE_Block2_start_1081_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1081_Update/$exit
      -- 
    ack_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_1, ack => convTranspose_CP_39_elements(306)); -- 
    req_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(306), ack => WPIPE_Block2_start_1084_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Update/req
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_update_start_
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_sample_completed_
      -- 
    ack_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_0, ack => convTranspose_CP_39_elements(307)); -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(307), ack => WPIPE_Block2_start_1084_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Sample/req
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1084_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_sample_start_
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_1, ack => convTranspose_CP_39_elements(308)); -- 
    req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => WPIPE_Block2_start_1087_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_update_start_
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Update/req
      -- 
    ack_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_0, ack => convTranspose_CP_39_elements(309)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => WPIPE_Block2_start_1087_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1087_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Sample/req
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_1, ack => convTranspose_CP_39_elements(310)); -- 
    req_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(310), ack => WPIPE_Block2_start_1090_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_update_start_
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Update/req
      -- 
    ack_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1090_inst_ack_0, ack => convTranspose_CP_39_elements(311)); -- 
    req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(311), ack => WPIPE_Block2_start_1090_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1090_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Sample/req
      -- 
    ack_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1090_inst_ack_1, ack => convTranspose_CP_39_elements(312)); -- 
    req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(312), ack => WPIPE_Block2_start_1093_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_update_start_
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Update/req
      -- 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1093_inst_ack_0, ack => convTranspose_CP_39_elements(313)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(313), ack => WPIPE_Block2_start_1093_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	317 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1093_Update/ack
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1093_inst_ack_1, ack => convTranspose_CP_39_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	469 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Sample/ra
      -- 
    ra_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_0, ack => convTranspose_CP_39_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	469 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Update/ca
      -- 
    ca_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_1, ack => convTranspose_CP_39_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	314 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Sample/req
      -- 
    req_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => WPIPE_Block2_start_1106_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(314) & convTranspose_CP_39_elements(316);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_update_start_
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Update/req
      -- 
    ack_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1106_inst_ack_0, ack => convTranspose_CP_39_elements(318)); -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(318), ack => WPIPE_Block2_start_1106_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1106_Update/ack
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1106_inst_ack_1, ack => convTranspose_CP_39_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	469 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Sample/ra
      -- 
    ra_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_0, ack => convTranspose_CP_39_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	469 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Update/ca
      -- 
    ca_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1111_inst_ack_1, ack => convTranspose_CP_39_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	319 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Sample/req
      -- 
    req_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(322), ack => WPIPE_Block2_start_1113_inst_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(319) & convTranspose_CP_39_elements(321);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_update_start_
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Update/req
      -- 
    ack_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1113_inst_ack_0, ack => convTranspose_CP_39_elements(323)); -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(323), ack => WPIPE_Block2_start_1113_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1113_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Sample/req
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1113_inst_ack_1, ack => convTranspose_CP_39_elements(324)); -- 
    req_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(324), ack => WPIPE_Block2_start_1116_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_update_start_
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Update/req
      -- 
    ack_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1116_inst_ack_0, ack => convTranspose_CP_39_elements(325)); -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(325), ack => WPIPE_Block2_start_1116_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1116_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Sample/req
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1116_inst_ack_1, ack => convTranspose_CP_39_elements(326)); -- 
    req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(326), ack => WPIPE_Block2_start_1119_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_update_start_
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Update/req
      -- 
    ack_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_0, ack => convTranspose_CP_39_elements(327)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(327), ack => WPIPE_Block2_start_1119_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1119_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Sample/req
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_1, ack => convTranspose_CP_39_elements(328)); -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(328), ack => WPIPE_Block2_start_1122_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_update_start_
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Update/req
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_0, ack => convTranspose_CP_39_elements(329)); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(329), ack => WPIPE_Block2_start_1122_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	373 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1122_Update/ack
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_1, ack => convTranspose_CP_39_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	469 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_update_start_
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Update/req
      -- 
    ack_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1125_inst_ack_0, ack => convTranspose_CP_39_elements(331)); -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(331), ack => WPIPE_Block3_start_1125_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Sample/req
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1125_inst_ack_1, ack => convTranspose_CP_39_elements(332)); -- 
    req_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(332), ack => WPIPE_Block3_start_1128_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_update_start_
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Update/req
      -- 
    ack_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1128_inst_ack_0, ack => convTranspose_CP_39_elements(333)); -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(333), ack => WPIPE_Block3_start_1128_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1128_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Sample/req
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1128_inst_ack_1, ack => convTranspose_CP_39_elements(334)); -- 
    req_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(334), ack => WPIPE_Block3_start_1131_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_update_start_
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Update/req
      -- 
    ack_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_0, ack => convTranspose_CP_39_elements(335)); -- 
    req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => WPIPE_Block3_start_1131_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1131_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Sample/req
      -- 
    ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_1, ack => convTranspose_CP_39_elements(336)); -- 
    req_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(336), ack => WPIPE_Block3_start_1134_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_update_start_
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Update/req
      -- 
    ack_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_0, ack => convTranspose_CP_39_elements(337)); -- 
    req_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(337), ack => WPIPE_Block3_start_1134_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1134_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Sample/req
      -- 
    ack_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_1, ack => convTranspose_CP_39_elements(338)); -- 
    req_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(338), ack => WPIPE_Block3_start_1137_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_update_start_
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Update/req
      -- 
    ack_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_0, ack => convTranspose_CP_39_elements(339)); -- 
    req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => WPIPE_Block3_start_1137_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1137_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Sample/req
      -- 
    ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_1, ack => convTranspose_CP_39_elements(340)); -- 
    req_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(340), ack => WPIPE_Block3_start_1140_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_update_start_
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Update/req
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_0, ack => convTranspose_CP_39_elements(341)); -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(341), ack => WPIPE_Block3_start_1140_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1140_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Sample/req
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_1, ack => convTranspose_CP_39_elements(342)); -- 
    req_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(342), ack => WPIPE_Block3_start_1143_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_update_start_
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Update/req
      -- 
    ack_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_0, ack => convTranspose_CP_39_elements(343)); -- 
    req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(343), ack => WPIPE_Block3_start_1143_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1143_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Sample/req
      -- 
    ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_1, ack => convTranspose_CP_39_elements(344)); -- 
    req_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(344), ack => WPIPE_Block3_start_1146_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_update_start_
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Update/req
      -- 
    ack_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1146_inst_ack_0, ack => convTranspose_CP_39_elements(345)); -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(345), ack => WPIPE_Block3_start_1146_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1146_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Sample/req
      -- 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1146_inst_ack_1, ack => convTranspose_CP_39_elements(346)); -- 
    req_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => WPIPE_Block3_start_1149_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_update_start_
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Update/req
      -- 
    ack_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1149_inst_ack_0, ack => convTranspose_CP_39_elements(347)); -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(347), ack => WPIPE_Block3_start_1149_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1149_Update/ack
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1149_inst_ack_1, ack => convTranspose_CP_39_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	469 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Sample/ra
      -- 
    ra_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1160_inst_ack_0, ack => convTranspose_CP_39_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	469 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Update/ca
      -- 
    ca_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1160_inst_ack_1, ack => convTranspose_CP_39_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Sample/req
      -- 
    req_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(351), ack => WPIPE_Block3_start_1162_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(348) & convTranspose_CP_39_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_update_start_
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Update/req
      -- 
    ack_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1162_inst_ack_0, ack => convTranspose_CP_39_elements(352)); -- 
    req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(352), ack => WPIPE_Block3_start_1162_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1162_Update/ack
      -- 
    ack_2682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1162_inst_ack_1, ack => convTranspose_CP_39_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	469 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Sample/ra
      -- 
    ra_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_0, ack => convTranspose_CP_39_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	469 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Update/ca
      -- 
    ca_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_1, ack => convTranspose_CP_39_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Sample/req
      -- 
    req_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(356), ack => WPIPE_Block3_start_1169_inst_req_0); -- 
    convTranspose_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(353) & convTranspose_CP_39_elements(355);
      gj_convTranspose_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_update_start_
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Sample/ack
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Update/req
      -- 
    ack_2705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1169_inst_ack_0, ack => convTranspose_CP_39_elements(357)); -- 
    req_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(357), ack => WPIPE_Block3_start_1169_inst_req_1); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1169_Update/ack
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Sample/req
      -- 
    ack_2710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1169_inst_ack_1, ack => convTranspose_CP_39_elements(358)); -- 
    req_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(358), ack => WPIPE_Block3_start_1172_inst_req_0); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_update_start_
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Update/req
      -- 
    ack_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1172_inst_ack_0, ack => convTranspose_CP_39_elements(359)); -- 
    req_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(359), ack => WPIPE_Block3_start_1172_inst_req_1); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1172_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Sample/req
      -- 
    ack_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1172_inst_ack_1, ack => convTranspose_CP_39_elements(360)); -- 
    req_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(360), ack => WPIPE_Block3_start_1175_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_update_start_
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Update/req
      -- 
    ack_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_0, ack => convTranspose_CP_39_elements(361)); -- 
    req_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(361), ack => WPIPE_Block3_start_1175_inst_req_1); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1175_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Sample/req
      -- 
    ack_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_1, ack => convTranspose_CP_39_elements(362)); -- 
    req_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(362), ack => WPIPE_Block3_start_1178_inst_req_0); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_update_start_
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Update/req
      -- 
    ack_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_0, ack => convTranspose_CP_39_elements(363)); -- 
    req_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(363), ack => WPIPE_Block3_start_1178_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	373 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1178_Update/ack
      -- 
    ack_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_1, ack => convTranspose_CP_39_elements(364)); -- 
    -- CP-element group 365:  transition  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	469 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_update_start_
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Sample/ra
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Update/cr
      -- 
    ra_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1182_inst_ack_0, ack => convTranspose_CP_39_elements(365)); -- 
    cr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(365), ack => RPIPE_Block0_done_1182_inst_req_1); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	373 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Update/ca
      -- 
    ca_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1182_inst_ack_1, ack => convTranspose_CP_39_elements(366)); -- 
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	469 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_update_start_
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Sample/ra
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Update/cr
      -- 
    ra_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1185_inst_ack_0, ack => convTranspose_CP_39_elements(367)); -- 
    cr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(367), ack => RPIPE_Block1_done_1185_inst_req_1); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	373 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Update/ca
      -- 
    ca_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1185_inst_ack_1, ack => convTranspose_CP_39_elements(368)); -- 
    -- CP-element group 369:  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	469 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_sample_completed_
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_update_start_
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Sample/ra
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Update/$entry
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Update/cr
      -- 
    ra_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1188_inst_ack_0, ack => convTranspose_CP_39_elements(369)); -- 
    cr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(369), ack => RPIPE_Block2_done_1188_inst_req_1); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	373 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_update_completed_
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Update/ca
      -- 
    ca_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1188_inst_ack_1, ack => convTranspose_CP_39_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	469 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_update_start_
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Sample/ra
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Update/$entry
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Update/cr
      -- 
    ra_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1191_inst_ack_0, ack => convTranspose_CP_39_elements(371)); -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(371), ack => RPIPE_Block3_done_1191_inst_req_1); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Update/ca
      -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1191_inst_ack_1, ack => convTranspose_CP_39_elements(372)); -- 
    -- CP-element group 373:  join  fork  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	364 
    -- CP-element group 373: 	366 
    -- CP-element group 373: 	368 
    -- CP-element group 373: 	370 
    -- CP-element group 373: 	372 
    -- CP-element group 373: 	234 
    -- CP-element group 373: 	262 
    -- CP-element group 373: 	296 
    -- CP-element group 373: 	330 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373: 	375 
    -- CP-element group 373: 	377 
    -- CP-element group 373: 	379 
    -- CP-element group 373: 	381 
    -- CP-element group 373: 	383 
    -- CP-element group 373: 	385 
    -- CP-element group 373:  members (25) 
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192__exit__
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251__entry__
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/$exit
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_Sample/crr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_Update/ccr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_Update/cr
      -- 
    crr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => call_stmt_1195_call_req_0); -- 
    ccr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => call_stmt_1195_call_req_1); -- 
    cr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1199_inst_req_1); -- 
    cr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1208_inst_req_1); -- 
    cr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1218_inst_req_1); -- 
    cr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1228_inst_req_1); -- 
    cr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => type_cast_1238_inst_req_1); -- 
    convTranspose_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(364) & convTranspose_CP_39_elements(366) & convTranspose_CP_39_elements(368) & convTranspose_CP_39_elements(370) & convTranspose_CP_39_elements(372) & convTranspose_CP_39_elements(234) & convTranspose_CP_39_elements(262) & convTranspose_CP_39_elements(296) & convTranspose_CP_39_elements(330);
      gj_convTranspose_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_Sample/$exit
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_Sample/cra
      -- 
    cra_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1195_call_ack_0, ack => convTranspose_CP_39_elements(374)); -- 
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/call_stmt_1195_Update/cca
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_Sample/rr
      -- 
    cca_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1195_call_ack_1, ack => convTranspose_CP_39_elements(375)); -- 
    rr_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(375), ack => type_cast_1199_inst_req_0); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_Sample/ra
      -- 
    ra_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1199_inst_ack_0, ack => convTranspose_CP_39_elements(376)); -- 
    -- CP-element group 377:  fork  transition  input  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	373 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377: 	380 
    -- CP-element group 377: 	382 
    -- CP-element group 377: 	384 
    -- CP-element group 377:  members (15) 
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1199_Update/ca
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_Sample/rr
      -- 
    ca_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1199_inst_ack_1, ack => convTranspose_CP_39_elements(377)); -- 
    rr_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1208_inst_req_0); -- 
    rr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1218_inst_req_0); -- 
    rr_2875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1228_inst_req_0); -- 
    rr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1238_inst_req_0); -- 
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_Sample/ra
      -- 
    ra_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1208_inst_ack_0, ack => convTranspose_CP_39_elements(378)); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	373 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	394 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1208_Update/ca
      -- 
    ca_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1208_inst_ack_1, ack => convTranspose_CP_39_elements(379)); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	377 
    -- CP-element group 380: successors 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_Sample/ra
      -- 
    ra_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1218_inst_ack_0, ack => convTranspose_CP_39_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	373 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	391 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1218_Update/ca
      -- 
    ca_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1218_inst_ack_1, ack => convTranspose_CP_39_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	377 
    -- CP-element group 382: successors 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_Sample/ra
      -- 
    ra_2876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1228_inst_ack_0, ack => convTranspose_CP_39_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	373 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	388 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1228_Update/ca
      -- 
    ca_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1228_inst_ack_1, ack => convTranspose_CP_39_elements(383)); -- 
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	377 
    -- CP-element group 384: successors 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_Sample/ra
      -- 
    ra_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => convTranspose_CP_39_elements(384)); -- 
    -- CP-element group 385:  transition  input  output  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	373 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (6) 
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/type_cast_1238_Update/ca
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_Sample/$entry
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_Sample/req
      -- 
    ca_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => convTranspose_CP_39_elements(385)); -- 
    req_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(385), ack => WPIPE_ConvTranspose_output_pipe_1240_inst_req_0); -- 
    -- CP-element group 386:  transition  input  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386:  members (6) 
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_Sample/ack
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_Update/req
      -- 
    ack_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1240_inst_ack_0, ack => convTranspose_CP_39_elements(386)); -- 
    req_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => WPIPE_ConvTranspose_output_pipe_1240_inst_req_1); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1240_Update/ack
      -- 
    ack_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1240_inst_ack_1, ack => convTranspose_CP_39_elements(387)); -- 
    -- CP-element group 388:  join  transition  output  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	383 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	389 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_sample_start_
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_Sample/$entry
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_Sample/req
      -- 
    req_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(388), ack => WPIPE_ConvTranspose_output_pipe_1243_inst_req_0); -- 
    convTranspose_cp_element_group_388: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_388"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(383) & convTranspose_CP_39_elements(387);
      gj_convTranspose_cp_element_group_388 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(388), clk => clk, reset => reset); --
    end block;
    -- CP-element group 389:  transition  input  output  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	388 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (6) 
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_sample_completed_
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_update_start_
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_Sample/ack
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_Update/$entry
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_Update/req
      -- 
    ack_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1243_inst_ack_0, ack => convTranspose_CP_39_elements(389)); -- 
    req_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => WPIPE_ConvTranspose_output_pipe_1243_inst_req_1); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_update_completed_
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1243_Update/ack
      -- 
    ack_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1243_inst_ack_1, ack => convTranspose_CP_39_elements(390)); -- 
    -- CP-element group 391:  join  transition  output  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	381 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_sample_start_
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_Sample/$entry
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_Sample/req
      -- 
    req_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(391), ack => WPIPE_ConvTranspose_output_pipe_1246_inst_req_0); -- 
    convTranspose_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(381) & convTranspose_CP_39_elements(390);
      gj_convTranspose_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  transition  input  output  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392:  members (6) 
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_update_start_
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_Sample/ack
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_Update/$entry
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_Update/req
      -- 
    ack_2932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1246_inst_ack_0, ack => convTranspose_CP_39_elements(392)); -- 
    req_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(392), ack => WPIPE_ConvTranspose_output_pipe_1246_inst_req_1); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	394 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1246_Update/ack
      -- 
    ack_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1246_inst_ack_1, ack => convTranspose_CP_39_elements(393)); -- 
    -- CP-element group 394:  join  transition  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	379 
    -- CP-element group 394: 	393 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_sample_start_
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_Sample/$entry
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_Sample/req
      -- 
    req_2945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(394), ack => WPIPE_ConvTranspose_output_pipe_1249_inst_req_0); -- 
    convTranspose_cp_element_group_394: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_394"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(379) & convTranspose_CP_39_elements(393);
      gj_convTranspose_cp_element_group_394 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(394), clk => clk, reset => reset); --
    end block;
    -- CP-element group 395:  transition  input  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (6) 
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_sample_completed_
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_update_start_
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_Sample/$exit
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_Sample/ack
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_Update/$entry
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_Update/req
      -- 
    ack_2946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1249_inst_ack_0, ack => convTranspose_CP_39_elements(395)); -- 
    req_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(395), ack => WPIPE_ConvTranspose_output_pipe_1249_inst_req_1); -- 
    -- CP-element group 396:  branch  transition  place  input  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396: 	398 
    -- CP-element group 396:  members (13) 
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251__exit__
      -- CP-element group 396: 	 branch_block_stmt_32/if_stmt_1253__entry__
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/$exit
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_update_completed_
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_Update/$exit
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_1195_to_assign_stmt_1251/WPIPE_ConvTranspose_output_pipe_1249_Update/ack
      -- CP-element group 396: 	 branch_block_stmt_32/if_stmt_1253_dead_link/$entry
      -- CP-element group 396: 	 branch_block_stmt_32/if_stmt_1253_eval_test/$entry
      -- CP-element group 396: 	 branch_block_stmt_32/if_stmt_1253_eval_test/$exit
      -- CP-element group 396: 	 branch_block_stmt_32/if_stmt_1253_eval_test/branch_req
      -- CP-element group 396: 	 branch_block_stmt_32/R_cmp264497_1254_place
      -- CP-element group 396: 	 branch_block_stmt_32/if_stmt_1253_if_link/$entry
      -- CP-element group 396: 	 branch_block_stmt_32/if_stmt_1253_else_link/$entry
      -- 
    ack_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1249_inst_ack_1, ack => convTranspose_CP_39_elements(396)); -- 
    branch_req_2959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(396), ack => if_stmt_1253_branch_req_0); -- 
    -- CP-element group 397:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	399 
    -- CP-element group 397: 	400 
    -- CP-element group 397:  members (18) 
      -- CP-element group 397: 	 branch_block_stmt_32/merge_stmt_1259__exit__
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294__entry__
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_update_start_
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_Update/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_Sample/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_Update/cr
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_sample_start_
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_Sample/rr
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/if_stmt_1253_if_link/$exit
      -- CP-element group 397: 	 branch_block_stmt_32/if_stmt_1253_if_link/if_choice_transition
      -- CP-element group 397: 	 branch_block_stmt_32/forx_xend273_bbx_xnph
      -- CP-element group 397: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 397: 	 branch_block_stmt_32/merge_stmt_1259_PhiReqMerge
      -- CP-element group 397: 	 branch_block_stmt_32/merge_stmt_1259_PhiAck/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/merge_stmt_1259_PhiAck/$exit
      -- CP-element group 397: 	 branch_block_stmt_32/merge_stmt_1259_PhiAck/dummy
      -- 
    if_choice_transition_2964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1253_branch_ack_1, ack => convTranspose_CP_39_elements(397)); -- 
    cr_2986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => type_cast_1280_inst_req_1); -- 
    rr_2981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => type_cast_1280_inst_req_0); -- 
    -- CP-element group 398:  transition  place  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	396 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	476 
    -- CP-element group 398:  members (5) 
      -- CP-element group 398: 	 branch_block_stmt_32/if_stmt_1253_else_link/$exit
      -- CP-element group 398: 	 branch_block_stmt_32/if_stmt_1253_else_link/else_choice_transition
      -- CP-element group 398: 	 branch_block_stmt_32/forx_xend273_forx_xend492
      -- CP-element group 398: 	 branch_block_stmt_32/forx_xend273_forx_xend492_PhiReq/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/forx_xend273_forx_xend492_PhiReq/$exit
      -- 
    else_choice_transition_2968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1253_branch_ack_0, ack => convTranspose_CP_39_elements(398)); -- 
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	397 
    -- CP-element group 399: successors 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_Sample/ra
      -- CP-element group 399: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_sample_completed_
      -- CP-element group 399: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_Sample/$exit
      -- 
    ra_2982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1280_inst_ack_0, ack => convTranspose_CP_39_elements(399)); -- 
    -- CP-element group 400:  transition  place  input  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	397 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	470 
    -- CP-element group 400:  members (9) 
      -- CP-element group 400: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294__exit__
      -- CP-element group 400: 	 branch_block_stmt_32/bbx_xnph_forx_xbody419
      -- CP-element group 400: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_update_completed_
      -- CP-element group 400: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_Update/$exit
      -- CP-element group 400: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/type_cast_1280_Update/ca
      -- CP-element group 400: 	 branch_block_stmt_32/assign_stmt_1265_to_assign_stmt_1294/$exit
      -- CP-element group 400: 	 branch_block_stmt_32/bbx_xnph_forx_xbody419_PhiReq/$entry
      -- CP-element group 400: 	 branch_block_stmt_32/bbx_xnph_forx_xbody419_PhiReq/phi_stmt_1297/$entry
      -- CP-element group 400: 	 branch_block_stmt_32/bbx_xnph_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/$entry
      -- 
    ca_2987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1280_inst_ack_1, ack => convTranspose_CP_39_elements(400)); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	475 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	446 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_final_index_sum_regn_Sample/ack
      -- CP-element group 401: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_final_index_sum_regn_Sample/$exit
      -- CP-element group 401: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_final_index_sum_regn_sample_complete
      -- 
    ack_3016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1309_index_offset_ack_0, ack => convTranspose_CP_39_elements(401)); -- 
    -- CP-element group 402:  transition  input  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	475 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (11) 
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_request/req
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_base_plus_offset/sum_rename_req
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_base_plus_offset/sum_rename_ack
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_request/$entry
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_final_index_sum_regn_Update/ack
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_base_plus_offset/$exit
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_base_plus_offset/$entry
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_final_index_sum_regn_Update/$exit
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_offset_calculated
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_root_address_calculated
      -- CP-element group 402: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_sample_start_
      -- 
    ack_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1309_index_offset_ack_1, ack => convTranspose_CP_39_elements(402)); -- 
    req_3030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(402), ack => addr_of_1310_final_reg_req_0); -- 
    -- CP-element group 403:  transition  input  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_request/ack
      -- CP-element group 403: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_request/$exit
      -- CP-element group 403: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_sample_completed_
      -- 
    ack_3031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1310_final_reg_ack_0, ack => convTranspose_CP_39_elements(403)); -- 
    -- CP-element group 404:  join  fork  transition  input  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	475 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (24) 
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_word_address_calculated
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_base_address_calculated
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_complete/$exit
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_complete/ack
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_sample_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Sample/word_access_start/word_0/rr
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Sample/word_access_start/word_0/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Sample/word_access_start/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Sample/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_word_addrgen/root_register_ack
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_word_addrgen/root_register_req
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_word_addrgen/$exit
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_update_completed_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_word_addrgen/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_base_plus_offset/sum_rename_ack
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_base_plus_offset/sum_rename_req
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_base_plus_offset/$exit
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_base_plus_offset/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_base_addr_resize/base_resize_ack
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_base_addr_resize/base_resize_req
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_base_addr_resize/$exit
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_base_addr_resize/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_base_address_resized
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_root_address_calculated
      -- 
    ack_3036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1310_final_reg_ack_1, ack => convTranspose_CP_39_elements(404)); -- 
    rr_3069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => ptr_deref_1314_load_0_req_0); -- 
    -- CP-element group 405:  transition  input  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405:  members (5) 
      -- CP-element group 405: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_sample_completed_
      -- CP-element group 405: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Sample/word_access_start/word_0/ra
      -- CP-element group 405: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Sample/word_access_start/word_0/$exit
      -- CP-element group 405: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Sample/word_access_start/$exit
      -- CP-element group 405: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Sample/$exit
      -- 
    ra_3070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1314_load_0_ack_0, ack => convTranspose_CP_39_elements(405)); -- 
    -- CP-element group 406:  fork  transition  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	475 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406: 	409 
    -- CP-element group 406: 	411 
    -- CP-element group 406: 	413 
    -- CP-element group 406: 	415 
    -- CP-element group 406: 	417 
    -- CP-element group 406: 	419 
    -- CP-element group 406: 	421 
    -- CP-element group 406:  members (33) 
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_sample_start_
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_update_completed_
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_sample_start_
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_sample_start_
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_sample_start_
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_sample_start_
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/ptr_deref_1314_Merge/merge_ack
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/ptr_deref_1314_Merge/merge_req
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/ptr_deref_1314_Merge/$exit
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/ptr_deref_1314_Merge/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/word_access_complete/word_0/ca
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_sample_start_
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/word_access_complete/word_0/$exit
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/word_access_complete/$exit
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/$exit
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_Sample/rr
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_sample_start_
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_Sample/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_sample_start_
      -- CP-element group 406: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_Sample/rr
      -- 
    ca_3081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1314_load_0_ack_1, ack => convTranspose_CP_39_elements(406)); -- 
    rr_3094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => type_cast_1318_inst_req_0); -- 
    rr_3108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => type_cast_1328_inst_req_0); -- 
    rr_3122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => type_cast_1338_inst_req_0); -- 
    rr_3136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => type_cast_1348_inst_req_0); -- 
    rr_3150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => type_cast_1358_inst_req_0); -- 
    rr_3164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => type_cast_1368_inst_req_0); -- 
    rr_3178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => type_cast_1378_inst_req_0); -- 
    rr_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => type_cast_1388_inst_req_0); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_Sample/ra
      -- CP-element group 407: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_Sample/$exit
      -- CP-element group 407: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_sample_completed_
      -- 
    ra_3095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1318_inst_ack_0, ack => convTranspose_CP_39_elements(407)); -- 
    -- CP-element group 408:  transition  input  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	475 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	443 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_Update/ca
      -- CP-element group 408: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_Update/$exit
      -- CP-element group 408: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_update_completed_
      -- 
    ca_3100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1318_inst_ack_1, ack => convTranspose_CP_39_elements(408)); -- 
    -- CP-element group 409:  transition  input  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	406 
    -- CP-element group 409: successors 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_Sample/ra
      -- CP-element group 409: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_Sample/$exit
      -- CP-element group 409: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_sample_completed_
      -- 
    ra_3109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1328_inst_ack_0, ack => convTranspose_CP_39_elements(409)); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	475 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	440 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_update_completed_
      -- CP-element group 410: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_Update/$exit
      -- CP-element group 410: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_Update/ca
      -- 
    ca_3114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1328_inst_ack_1, ack => convTranspose_CP_39_elements(410)); -- 
    -- CP-element group 411:  transition  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	406 
    -- CP-element group 411: successors 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_Sample/$exit
      -- CP-element group 411: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_sample_completed_
      -- CP-element group 411: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_Sample/ra
      -- 
    ra_3123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_0, ack => convTranspose_CP_39_elements(411)); -- 
    -- CP-element group 412:  transition  input  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	475 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	437 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_update_completed_
      -- CP-element group 412: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_Update/ca
      -- CP-element group 412: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_Update/$exit
      -- 
    ca_3128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_1, ack => convTranspose_CP_39_elements(412)); -- 
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	406 
    -- CP-element group 413: successors 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_Sample/ra
      -- CP-element group 413: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_Sample/$exit
      -- CP-element group 413: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_sample_completed_
      -- 
    ra_3137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1348_inst_ack_0, ack => convTranspose_CP_39_elements(413)); -- 
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	475 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	434 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_Update/ca
      -- CP-element group 414: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_Update/$exit
      -- CP-element group 414: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_update_completed_
      -- 
    ca_3142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1348_inst_ack_1, ack => convTranspose_CP_39_elements(414)); -- 
    -- CP-element group 415:  transition  input  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	406 
    -- CP-element group 415: successors 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_Sample/ra
      -- CP-element group 415: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_Sample/$exit
      -- CP-element group 415: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_sample_completed_
      -- 
    ra_3151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_0, ack => convTranspose_CP_39_elements(415)); -- 
    -- CP-element group 416:  transition  input  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	475 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	431 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_Update/ca
      -- CP-element group 416: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_update_completed_
      -- 
    ca_3156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_1, ack => convTranspose_CP_39_elements(416)); -- 
    -- CP-element group 417:  transition  input  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	406 
    -- CP-element group 417: successors 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_Sample/ra
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_Sample/$exit
      -- CP-element group 417: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_sample_completed_
      -- 
    ra_3165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_0, ack => convTranspose_CP_39_elements(417)); -- 
    -- CP-element group 418:  transition  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	475 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	428 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_Update/ca
      -- CP-element group 418: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_Update/$exit
      -- CP-element group 418: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_update_completed_
      -- 
    ca_3170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_1, ack => convTranspose_CP_39_elements(418)); -- 
    -- CP-element group 419:  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	406 
    -- CP-element group 419: successors 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_Sample/ra
      -- CP-element group 419: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_sample_completed_
      -- 
    ra_3179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_0, ack => convTranspose_CP_39_elements(419)); -- 
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	475 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	425 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_update_completed_
      -- CP-element group 420: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_Update/ca
      -- 
    ca_3184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_1, ack => convTranspose_CP_39_elements(420)); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	406 
    -- CP-element group 421: successors 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_Sample/ra
      -- CP-element group 421: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_Sample/$exit
      -- CP-element group 421: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_sample_completed_
      -- 
    ra_3193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_0, ack => convTranspose_CP_39_elements(421)); -- 
    -- CP-element group 422:  transition  input  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	475 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (6) 
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_Sample/req
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_Sample/$entry
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_sample_start_
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_Update/ca
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_Update/$exit
      -- CP-element group 422: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_update_completed_
      -- 
    ca_3198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_1, ack => convTranspose_CP_39_elements(422)); -- 
    req_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(422), ack => WPIPE_ConvTranspose_output_pipe_1390_inst_req_0); -- 
    -- CP-element group 423:  transition  input  output  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (6) 
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_Update/req
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_Update/$entry
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_Sample/ack
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_Sample/$exit
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_update_start_
      -- CP-element group 423: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_sample_completed_
      -- 
    ack_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1390_inst_ack_0, ack => convTranspose_CP_39_elements(423)); -- 
    req_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(423), ack => WPIPE_ConvTranspose_output_pipe_1390_inst_req_1); -- 
    -- CP-element group 424:  transition  input  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_Update/ack
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_Update/$exit
      -- CP-element group 424: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1390_update_completed_
      -- 
    ack_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1390_inst_ack_1, ack => convTranspose_CP_39_elements(424)); -- 
    -- CP-element group 425:  join  transition  output  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	420 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_Sample/$entry
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_Sample/req
      -- CP-element group 425: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_sample_start_
      -- 
    req_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(425), ack => WPIPE_ConvTranspose_output_pipe_1393_inst_req_0); -- 
    convTranspose_cp_element_group_425: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_425"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(420) & convTranspose_CP_39_elements(424);
      gj_convTranspose_cp_element_group_425 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(425), clk => clk, reset => reset); --
    end block;
    -- CP-element group 426:  transition  input  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426:  members (6) 
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_Sample/$exit
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_update_start_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_Sample/ack
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_sample_completed_
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_Update/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_Update/req
      -- 
    ack_3221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1393_inst_ack_0, ack => convTranspose_CP_39_elements(426)); -- 
    req_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => WPIPE_ConvTranspose_output_pipe_1393_inst_req_1); -- 
    -- CP-element group 427:  transition  input  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_update_completed_
      -- CP-element group 427: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_Update/ack
      -- CP-element group 427: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1393_Update/$exit
      -- 
    ack_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1393_inst_ack_1, ack => convTranspose_CP_39_elements(427)); -- 
    -- CP-element group 428:  join  transition  output  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	418 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_Sample/req
      -- CP-element group 428: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_Sample/$entry
      -- CP-element group 428: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_sample_start_
      -- 
    req_3234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(428), ack => WPIPE_ConvTranspose_output_pipe_1396_inst_req_0); -- 
    convTranspose_cp_element_group_428: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_428"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(418) & convTranspose_CP_39_elements(427);
      gj_convTranspose_cp_element_group_428 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(428), clk => clk, reset => reset); --
    end block;
    -- CP-element group 429:  transition  input  output  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	428 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429:  members (6) 
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_Update/req
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_Sample/ack
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_Update/$entry
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_Sample/$exit
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_update_start_
      -- CP-element group 429: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_sample_completed_
      -- 
    ack_3235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1396_inst_ack_0, ack => convTranspose_CP_39_elements(429)); -- 
    req_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => WPIPE_ConvTranspose_output_pipe_1396_inst_req_1); -- 
    -- CP-element group 430:  transition  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	431 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_Update/ack
      -- CP-element group 430: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_Update/$exit
      -- CP-element group 430: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1396_update_completed_
      -- 
    ack_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1396_inst_ack_1, ack => convTranspose_CP_39_elements(430)); -- 
    -- CP-element group 431:  join  transition  output  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	416 
    -- CP-element group 431: 	430 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	432 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_sample_start_
      -- CP-element group 431: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_Sample/req
      -- CP-element group 431: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_Sample/$entry
      -- 
    req_3248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(431), ack => WPIPE_ConvTranspose_output_pipe_1399_inst_req_0); -- 
    convTranspose_cp_element_group_431: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_431"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(416) & convTranspose_CP_39_elements(430);
      gj_convTranspose_cp_element_group_431 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(431), clk => clk, reset => reset); --
    end block;
    -- CP-element group 432:  transition  input  output  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	431 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	433 
    -- CP-element group 432:  members (6) 
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_sample_completed_
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_update_start_
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_Update/req
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_Update/$entry
      -- CP-element group 432: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_Sample/ack
      -- 
    ack_3249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1399_inst_ack_0, ack => convTranspose_CP_39_elements(432)); -- 
    req_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(432), ack => WPIPE_ConvTranspose_output_pipe_1399_inst_req_1); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	432 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	434 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_update_completed_
      -- CP-element group 433: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_Update/ack
      -- CP-element group 433: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1399_Update/$exit
      -- 
    ack_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1399_inst_ack_1, ack => convTranspose_CP_39_elements(433)); -- 
    -- CP-element group 434:  join  transition  output  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	414 
    -- CP-element group 434: 	433 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	435 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_Sample/$entry
      -- CP-element group 434: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_Sample/req
      -- CP-element group 434: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_sample_start_
      -- 
    req_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(434), ack => WPIPE_ConvTranspose_output_pipe_1402_inst_req_0); -- 
    convTranspose_cp_element_group_434: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_434"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(414) & convTranspose_CP_39_elements(433);
      gj_convTranspose_cp_element_group_434 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(434), clk => clk, reset => reset); --
    end block;
    -- CP-element group 435:  transition  input  output  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	434 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435:  members (6) 
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_Sample/$exit
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_Sample/ack
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_Update/$entry
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_update_start_
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_sample_completed_
      -- CP-element group 435: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_Update/req
      -- 
    ack_3263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1402_inst_ack_0, ack => convTranspose_CP_39_elements(435)); -- 
    req_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(435), ack => WPIPE_ConvTranspose_output_pipe_1402_inst_req_1); -- 
    -- CP-element group 436:  transition  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	435 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	437 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_update_completed_
      -- CP-element group 436: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_Update/ack
      -- CP-element group 436: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1402_Update/$exit
      -- 
    ack_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1402_inst_ack_1, ack => convTranspose_CP_39_elements(436)); -- 
    -- CP-element group 437:  join  transition  output  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	412 
    -- CP-element group 437: 	436 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	438 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_Sample/req
      -- CP-element group 437: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_Sample/$entry
      -- CP-element group 437: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_sample_start_
      -- 
    req_3276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(437), ack => WPIPE_ConvTranspose_output_pipe_1405_inst_req_0); -- 
    convTranspose_cp_element_group_437: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_437"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(412) & convTranspose_CP_39_elements(436);
      gj_convTranspose_cp_element_group_437 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(437), clk => clk, reset => reset); --
    end block;
    -- CP-element group 438:  transition  input  output  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	437 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	439 
    -- CP-element group 438:  members (6) 
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_Update/req
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_Sample/ack
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_Sample/$exit
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_update_start_
      -- CP-element group 438: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_sample_completed_
      -- 
    ack_3277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1405_inst_ack_0, ack => convTranspose_CP_39_elements(438)); -- 
    req_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => WPIPE_ConvTranspose_output_pipe_1405_inst_req_1); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	438 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	440 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_Update/ack
      -- CP-element group 439: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_Update/$exit
      -- CP-element group 439: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1405_update_completed_
      -- 
    ack_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1405_inst_ack_1, ack => convTranspose_CP_39_elements(439)); -- 
    -- CP-element group 440:  join  transition  output  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	410 
    -- CP-element group 440: 	439 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	441 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_Sample/req
      -- CP-element group 440: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_Sample/$entry
      -- CP-element group 440: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_sample_start_
      -- 
    req_3290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(440), ack => WPIPE_ConvTranspose_output_pipe_1408_inst_req_0); -- 
    convTranspose_cp_element_group_440: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_440"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(410) & convTranspose_CP_39_elements(439);
      gj_convTranspose_cp_element_group_440 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(440), clk => clk, reset => reset); --
    end block;
    -- CP-element group 441:  transition  input  output  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	440 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	442 
    -- CP-element group 441:  members (6) 
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_Update/req
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_Update/$entry
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_Sample/ack
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_Sample/$exit
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_update_start_
      -- CP-element group 441: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_sample_completed_
      -- 
    ack_3291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1408_inst_ack_0, ack => convTranspose_CP_39_elements(441)); -- 
    req_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(441), ack => WPIPE_ConvTranspose_output_pipe_1408_inst_req_1); -- 
    -- CP-element group 442:  transition  input  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	441 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	443 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_Update/ack
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_Update/$exit
      -- CP-element group 442: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1408_update_completed_
      -- 
    ack_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1408_inst_ack_1, ack => convTranspose_CP_39_elements(442)); -- 
    -- CP-element group 443:  join  transition  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	408 
    -- CP-element group 443: 	442 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	444 
    -- CP-element group 443:  members (3) 
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_Sample/req
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_Sample/$entry
      -- CP-element group 443: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_sample_start_
      -- 
    req_3304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(443), ack => WPIPE_ConvTranspose_output_pipe_1411_inst_req_0); -- 
    convTranspose_cp_element_group_443: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_443"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(408) & convTranspose_CP_39_elements(442);
      gj_convTranspose_cp_element_group_443 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(443), clk => clk, reset => reset); --
    end block;
    -- CP-element group 444:  transition  input  output  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	443 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	445 
    -- CP-element group 444:  members (6) 
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_Update/req
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_Update/$entry
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_Sample/ack
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_Sample/$exit
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_update_start_
      -- CP-element group 444: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_sample_completed_
      -- 
    ack_3305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1411_inst_ack_0, ack => convTranspose_CP_39_elements(444)); -- 
    req_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(444), ack => WPIPE_ConvTranspose_output_pipe_1411_inst_req_1); -- 
    -- CP-element group 445:  transition  input  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	444 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_Update/ack
      -- CP-element group 445: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_Update/$exit
      -- CP-element group 445: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/WPIPE_ConvTranspose_output_pipe_1411_update_completed_
      -- 
    ack_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1411_inst_ack_1, ack => convTranspose_CP_39_elements(445)); -- 
    -- CP-element group 446:  branch  join  transition  place  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	401 
    -- CP-element group 446: 	445 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446: 	448 
    -- CP-element group 446:  members (10) 
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424__exit__
      -- CP-element group 446: 	 branch_block_stmt_32/if_stmt_1425__entry__
      -- CP-element group 446: 	 branch_block_stmt_32/R_exitcond1_1426_place
      -- CP-element group 446: 	 branch_block_stmt_32/if_stmt_1425_else_link/$entry
      -- CP-element group 446: 	 branch_block_stmt_32/if_stmt_1425_if_link/$entry
      -- CP-element group 446: 	 branch_block_stmt_32/if_stmt_1425_eval_test/branch_req
      -- CP-element group 446: 	 branch_block_stmt_32/if_stmt_1425_eval_test/$exit
      -- CP-element group 446: 	 branch_block_stmt_32/if_stmt_1425_eval_test/$entry
      -- CP-element group 446: 	 branch_block_stmt_32/if_stmt_1425_dead_link/$entry
      -- CP-element group 446: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/$exit
      -- 
    branch_req_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(446), ack => if_stmt_1425_branch_req_0); -- 
    convTranspose_cp_element_group_446: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_446"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(401) & convTranspose_CP_39_elements(445);
      gj_convTranspose_cp_element_group_446 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(446), clk => clk, reset => reset); --
    end block;
    -- CP-element group 447:  merge  transition  place  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	476 
    -- CP-element group 447:  members (13) 
      -- CP-element group 447: 	 branch_block_stmt_32/merge_stmt_1431__exit__
      -- CP-element group 447: 	 branch_block_stmt_32/forx_xend492x_xloopexit_forx_xend492
      -- CP-element group 447: 	 branch_block_stmt_32/forx_xbody419_forx_xend492x_xloopexit
      -- CP-element group 447: 	 branch_block_stmt_32/if_stmt_1425_if_link/if_choice_transition
      -- CP-element group 447: 	 branch_block_stmt_32/if_stmt_1425_if_link/$exit
      -- CP-element group 447: 	 branch_block_stmt_32/forx_xbody419_forx_xend492x_xloopexit_PhiReq/$entry
      -- CP-element group 447: 	 branch_block_stmt_32/forx_xbody419_forx_xend492x_xloopexit_PhiReq/$exit
      -- CP-element group 447: 	 branch_block_stmt_32/merge_stmt_1431_PhiReqMerge
      -- CP-element group 447: 	 branch_block_stmt_32/merge_stmt_1431_PhiAck/$entry
      -- CP-element group 447: 	 branch_block_stmt_32/merge_stmt_1431_PhiAck/$exit
      -- CP-element group 447: 	 branch_block_stmt_32/merge_stmt_1431_PhiAck/dummy
      -- CP-element group 447: 	 branch_block_stmt_32/forx_xend492x_xloopexit_forx_xend492_PhiReq/$entry
      -- CP-element group 447: 	 branch_block_stmt_32/forx_xend492x_xloopexit_forx_xend492_PhiReq/$exit
      -- 
    if_choice_transition_3323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1425_branch_ack_1, ack => convTranspose_CP_39_elements(447)); -- 
    -- CP-element group 448:  fork  transition  place  input  output  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	446 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	471 
    -- CP-element group 448: 	472 
    -- CP-element group 448:  members (12) 
      -- CP-element group 448: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419
      -- CP-element group 448: 	 branch_block_stmt_32/if_stmt_1425_else_link/else_choice_transition
      -- CP-element group 448: 	 branch_block_stmt_32/if_stmt_1425_else_link/$exit
      -- CP-element group 448: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/$entry
      -- CP-element group 448: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/$entry
      -- CP-element group 448: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/$entry
      -- CP-element group 448: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/$entry
      -- CP-element group 448: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/$entry
      -- CP-element group 448: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Sample/$entry
      -- CP-element group 448: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Sample/rr
      -- CP-element group 448: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Update/$entry
      -- CP-element group 448: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1425_branch_ack_0, ack => convTranspose_CP_39_elements(448)); -- 
    rr_3602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(448), ack => type_cast_1303_inst_req_0); -- 
    cr_3607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(448), ack => type_cast_1303_inst_req_1); -- 
    -- CP-element group 449:  merge  branch  transition  place  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	165 
    -- CP-element group 449: 	120 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	121 
    -- CP-element group 449: 	122 
    -- CP-element group 449:  members (17) 
      -- CP-element group 449: 	 branch_block_stmt_32/merge_stmt_424__exit__
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_430__entry__
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_430__exit__
      -- CP-element group 449: 	 branch_block_stmt_32/if_stmt_431__entry__
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_430/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/assign_stmt_430/$exit
      -- CP-element group 449: 	 branch_block_stmt_32/if_stmt_431_dead_link/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/if_stmt_431_eval_test/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/if_stmt_431_eval_test/$exit
      -- CP-element group 449: 	 branch_block_stmt_32/if_stmt_431_eval_test/branch_req
      -- CP-element group 449: 	 branch_block_stmt_32/R_cmp194501_432_place
      -- CP-element group 449: 	 branch_block_stmt_32/if_stmt_431_if_link/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/if_stmt_431_else_link/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/merge_stmt_424_PhiAck/dummy
      -- CP-element group 449: 	 branch_block_stmt_32/merge_stmt_424_PhiAck/$exit
      -- CP-element group 449: 	 branch_block_stmt_32/merge_stmt_424_PhiAck/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/merge_stmt_424_PhiReqMerge
      -- 
    branch_req_925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(449), ack => if_stmt_431_branch_req_0); -- 
    convTranspose_CP_39_elements(449) <= OrReduce(convTranspose_CP_39_elements(165) & convTranspose_CP_39_elements(120));
    -- CP-element group 450:  transition  output  delay-element  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	124 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	454 
    -- CP-element group 450:  members (5) 
      -- CP-element group 450: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_req
      -- CP-element group 450: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_473_konst_delay_trans
      -- CP-element group 450: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$exit
      -- CP-element group 450: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody_PhiReq/phi_stmt_469/$exit
      -- CP-element group 450: 	 branch_block_stmt_32/bbx_xnph507_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_469_req_3375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_469_req_3375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(450), ack => phi_stmt_469_req_0); -- 
    -- Element group convTranspose_CP_39_elements(450) is a control-delay.
    cp_element_450_delay: control_delay_element  generic map(name => " 450_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(124), ack => convTranspose_CP_39_elements(450), clk => clk, reset =>reset);
    -- CP-element group 451:  transition  input  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	166 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	453 
    -- CP-element group 451:  members (2) 
      -- CP-element group 451: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/$exit
      -- CP-element group 451: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Sample/ra
      -- 
    ra_3395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_475_inst_ack_0, ack => convTranspose_CP_39_elements(451)); -- 
    -- CP-element group 452:  transition  input  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	166 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (2) 
      -- CP-element group 452: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/$exit
      -- CP-element group 452: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/Update/ca
      -- 
    ca_3400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_475_inst_ack_1, ack => convTranspose_CP_39_elements(452)); -- 
    -- CP-element group 453:  join  transition  output  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	451 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (6) 
      -- CP-element group 453: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 453: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/$exit
      -- CP-element group 453: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/$exit
      -- CP-element group 453: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/$exit
      -- CP-element group 453: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_sources/type_cast_475/SplitProtocol/$exit
      -- CP-element group 453: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_469/phi_stmt_469_req
      -- 
    phi_stmt_469_req_3401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_469_req_3401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(453), ack => phi_stmt_469_req_1); -- 
    convTranspose_cp_element_group_453: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_453"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(451) & convTranspose_CP_39_elements(452);
      gj_convTranspose_cp_element_group_453 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(453), clk => clk, reset => reset); --
    end block;
    -- CP-element group 454:  merge  transition  place  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	450 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (2) 
      -- CP-element group 454: 	 branch_block_stmt_32/merge_stmt_468_PhiReqMerge
      -- CP-element group 454: 	 branch_block_stmt_32/merge_stmt_468_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(454) <= OrReduce(convTranspose_CP_39_elements(450) & convTranspose_CP_39_elements(453));
    -- CP-element group 455:  fork  transition  place  input  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	163 
    -- CP-element group 455: 	125 
    -- CP-element group 455: 	126 
    -- CP-element group 455: 	128 
    -- CP-element group 455: 	129 
    -- CP-element group 455: 	132 
    -- CP-element group 455: 	136 
    -- CP-element group 455: 	140 
    -- CP-element group 455: 	144 
    -- CP-element group 455: 	148 
    -- CP-element group 455: 	152 
    -- CP-element group 455: 	156 
    -- CP-element group 455: 	160 
    -- CP-element group 455:  members (56) 
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/merge_stmt_468__exit__
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631__entry__
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/cr
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_538_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/cr
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/word_0/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/word_access_complete/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/cr
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/ptr_deref_618_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/cr
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_574_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_610_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/cr
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_556_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_592_Update/cr
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resized_1
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scaled_1
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_computed_1
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/$exit
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/index_resize_req
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_resize_1/index_resize_ack
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/$exit
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/scale_rename_req
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_index_scale_1/scale_rename_ack
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_update_start
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Sample/req
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/array_obj_ref_481_final_index_sum_regn_Update/req
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/addr_of_482_complete/req
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_sample_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/RPIPE_ConvTranspose_input_pipe_485_Sample/rr
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_489_Update/cr
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_502_Update/cr
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_update_start_
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/assign_stmt_483_to_assign_stmt_631/type_cast_520_Update/cr
      -- CP-element group 455: 	 branch_block_stmt_32/merge_stmt_468_PhiAck/$exit
      -- CP-element group 455: 	 branch_block_stmt_32/merge_stmt_468_PhiAck/phi_stmt_469_ack
      -- 
    phi_stmt_469_ack_3406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_469_ack_0, ack => convTranspose_CP_39_elements(455)); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => type_cast_538_inst_req_1); -- 
    cr_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => ptr_deref_618_store_0_req_1); -- 
    cr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => type_cast_610_inst_req_1); -- 
    cr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => type_cast_574_inst_req_1); -- 
    cr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => type_cast_556_inst_req_1); -- 
    cr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => type_cast_592_inst_req_1); -- 
    req_981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => array_obj_ref_481_index_offset_req_0); -- 
    req_986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => array_obj_ref_481_index_offset_req_1); -- 
    req_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => addr_of_482_final_reg_req_1); -- 
    rr_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => RPIPE_ConvTranspose_input_pipe_485_inst_req_0); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => type_cast_489_inst_req_1); -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => type_cast_502_inst_req_1); -- 
    cr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => type_cast_520_inst_req_1); -- 
    -- CP-element group 456:  transition  output  delay-element  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	168 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	460 
    -- CP-element group 456:  members (5) 
      -- CP-element group 456: 	 branch_block_stmt_32/bbx_xnph503_forx_xbody196_PhiReq/$exit
      -- CP-element group 456: 	 branch_block_stmt_32/bbx_xnph503_forx_xbody196_PhiReq/phi_stmt_676/$exit
      -- CP-element group 456: 	 branch_block_stmt_32/bbx_xnph503_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$exit
      -- CP-element group 456: 	 branch_block_stmt_32/bbx_xnph503_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_682_konst_delay_trans
      -- CP-element group 456: 	 branch_block_stmt_32/bbx_xnph503_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_req
      -- 
    phi_stmt_676_req_3429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_676_req_3429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(456), ack => phi_stmt_676_req_1); -- 
    -- Element group convTranspose_CP_39_elements(456) is a control-delay.
    cp_element_456_delay: control_delay_element  generic map(name => " 456_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(168), ack => convTranspose_CP_39_elements(456), clk => clk, reset =>reset);
    -- CP-element group 457:  transition  input  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	210 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	459 
    -- CP-element group 457:  members (2) 
      -- CP-element group 457: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/$exit
      -- CP-element group 457: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Sample/ra
      -- 
    ra_3449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_0, ack => convTranspose_CP_39_elements(457)); -- 
    -- CP-element group 458:  transition  input  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	210 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458:  members (2) 
      -- CP-element group 458: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/$exit
      -- CP-element group 458: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/Update/ca
      -- 
    ca_3454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_1, ack => convTranspose_CP_39_elements(458)); -- 
    -- CP-element group 459:  join  transition  output  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	457 
    -- CP-element group 459: 	458 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	460 
    -- CP-element group 459:  members (6) 
      -- CP-element group 459: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 459: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/$exit
      -- CP-element group 459: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/$exit
      -- CP-element group 459: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/$exit
      -- CP-element group 459: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_sources/type_cast_679/SplitProtocol/$exit
      -- CP-element group 459: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_676/phi_stmt_676_req
      -- 
    phi_stmt_676_req_3455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_676_req_3455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(459), ack => phi_stmt_676_req_0); -- 
    convTranspose_cp_element_group_459: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_459"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(457) & convTranspose_CP_39_elements(458);
      gj_convTranspose_cp_element_group_459 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(459), clk => clk, reset => reset); --
    end block;
    -- CP-element group 460:  merge  transition  place  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	456 
    -- CP-element group 460: 	459 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460:  members (2) 
      -- CP-element group 460: 	 branch_block_stmt_32/merge_stmt_675_PhiReqMerge
      -- CP-element group 460: 	 branch_block_stmt_32/merge_stmt_675_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(460) <= OrReduce(convTranspose_CP_39_elements(456) & convTranspose_CP_39_elements(459));
    -- CP-element group 461:  fork  transition  place  input  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	196 
    -- CP-element group 461: 	200 
    -- CP-element group 461: 	204 
    -- CP-element group 461: 	207 
    -- CP-element group 461: 	192 
    -- CP-element group 461: 	169 
    -- CP-element group 461: 	170 
    -- CP-element group 461: 	172 
    -- CP-element group 461: 	173 
    -- CP-element group 461: 	176 
    -- CP-element group 461: 	180 
    -- CP-element group 461: 	184 
    -- CP-element group 461: 	188 
    -- CP-element group 461:  members (56) 
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/cr
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/merge_stmt_675__exit__
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838__entry__
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/cr
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resized_1
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/req
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_709_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/rr
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_complete/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/addr_of_689_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/req
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_sample_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/RPIPE_ConvTranspose_input_pipe_692_Sample/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/cr
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/req
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_727_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_Sample/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_final_index_sum_regn_update_start
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/scale_rename_ack
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/scale_rename_req
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/$exit
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scale_1/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/index_resize_ack
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/index_resize_req
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_696_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/$exit
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_resize_1/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_computed_1
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/array_obj_ref_688_index_scaled_1
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_745_Update/cr
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_763_Update/cr
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_781_Update/cr
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_799_Update/cr
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/type_cast_817_Update/cr
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_update_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_690_to_assign_stmt_838/ptr_deref_825_Update/word_access_complete/word_0/cr
      -- CP-element group 461: 	 branch_block_stmt_32/merge_stmt_675_PhiAck/$exit
      -- CP-element group 461: 	 branch_block_stmt_32/merge_stmt_675_PhiAck/phi_stmt_676_ack
      -- 
    phi_stmt_676_ack_3460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_676_ack_0, ack => convTranspose_CP_39_elements(461)); -- 
    cr_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => type_cast_727_inst_req_1); -- 
    cr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => type_cast_709_inst_req_1); -- 
    req_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => addr_of_689_final_reg_req_1); -- 
    rr_1369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => RPIPE_ConvTranspose_input_pipe_692_inst_req_0); -- 
    req_1345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => array_obj_ref_688_index_offset_req_1); -- 
    cr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => type_cast_696_inst_req_1); -- 
    req_1340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => array_obj_ref_688_index_offset_req_0); -- 
    cr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => type_cast_745_inst_req_1); -- 
    cr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => type_cast_763_inst_req_1); -- 
    cr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => type_cast_781_inst_req_1); -- 
    cr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => type_cast_799_inst_req_1); -- 
    cr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => type_cast_817_inst_req_1); -- 
    cr_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => ptr_deref_825_store_0_req_1); -- 
    -- CP-element group 462:  merge  fork  transition  place  output  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	209 
    -- CP-element group 462: 	122 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	211 
    -- CP-element group 462: 	212 
    -- CP-element group 462: 	213 
    -- CP-element group 462: 	214 
    -- CP-element group 462: 	215 
    -- CP-element group 462: 	216 
    -- CP-element group 462:  members (25) 
      -- CP-element group 462: 	 branch_block_stmt_32/merge_stmt_847__exit__
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875__entry__
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/$entry
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_sample_start_
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_update_start_
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/$entry
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Sample/rr
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/$entry
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_850_Update/cr
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_sample_start_
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_update_start_
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/$entry
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Sample/rr
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/$entry
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_854_Update/cr
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_sample_start_
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_update_start_
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/$entry
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Sample/rr
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/$entry
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_851_to_assign_stmt_875/type_cast_858_Update/cr
      -- CP-element group 462: 	 branch_block_stmt_32/merge_stmt_847_PhiReqMerge
      -- CP-element group 462: 	 branch_block_stmt_32/merge_stmt_847_PhiAck/$entry
      -- CP-element group 462: 	 branch_block_stmt_32/merge_stmt_847_PhiAck/$exit
      -- CP-element group 462: 	 branch_block_stmt_32/merge_stmt_847_PhiAck/dummy
      -- 
    rr_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(462), ack => type_cast_850_inst_req_0); -- 
    cr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(462), ack => type_cast_850_inst_req_1); -- 
    rr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(462), ack => type_cast_854_inst_req_0); -- 
    cr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(462), ack => type_cast_854_inst_req_1); -- 
    rr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(462), ack => type_cast_858_inst_req_0); -- 
    cr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(462), ack => type_cast_858_inst_req_1); -- 
    convTranspose_CP_39_elements(462) <= OrReduce(convTranspose_CP_39_elements(209) & convTranspose_CP_39_elements(122));
    -- CP-element group 463:  transition  output  delay-element  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	221 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	467 
    -- CP-element group 463:  members (5) 
      -- CP-element group 463: 	 branch_block_stmt_32/bbx_xnph499_forx_xbody266_PhiReq/$exit
      -- CP-element group 463: 	 branch_block_stmt_32/bbx_xnph499_forx_xbody266_PhiReq/phi_stmt_920/$exit
      -- CP-element group 463: 	 branch_block_stmt_32/bbx_xnph499_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$exit
      -- CP-element group 463: 	 branch_block_stmt_32/bbx_xnph499_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_926_konst_delay_trans
      -- CP-element group 463: 	 branch_block_stmt_32/bbx_xnph499_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_req
      -- 
    phi_stmt_920_req_3506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_920_req_3506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(463), ack => phi_stmt_920_req_1); -- 
    -- Element group convTranspose_CP_39_elements(463) is a control-delay.
    cp_element_463_delay: control_delay_element  generic map(name => " 463_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(221), ack => convTranspose_CP_39_elements(463), clk => clk, reset =>reset);
    -- CP-element group 464:  transition  input  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	230 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	466 
    -- CP-element group 464:  members (2) 
      -- CP-element group 464: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/$exit
      -- CP-element group 464: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Sample/ra
      -- 
    ra_3526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_0, ack => convTranspose_CP_39_elements(464)); -- 
    -- CP-element group 465:  transition  input  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	230 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	466 
    -- CP-element group 465:  members (2) 
      -- CP-element group 465: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/$exit
      -- CP-element group 465: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/Update/ca
      -- 
    ca_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_1, ack => convTranspose_CP_39_elements(465)); -- 
    -- CP-element group 466:  join  transition  output  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	464 
    -- CP-element group 466: 	465 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	467 
    -- CP-element group 466:  members (6) 
      -- CP-element group 466: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 466: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/$exit
      -- CP-element group 466: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/$exit
      -- CP-element group 466: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/$exit
      -- CP-element group 466: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_sources/type_cast_923/SplitProtocol/$exit
      -- CP-element group 466: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_920/phi_stmt_920_req
      -- 
    phi_stmt_920_req_3532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_920_req_3532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(466), ack => phi_stmt_920_req_0); -- 
    convTranspose_cp_element_group_466: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_466"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(464) & convTranspose_CP_39_elements(465);
      gj_convTranspose_cp_element_group_466 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(466), clk => clk, reset => reset); --
    end block;
    -- CP-element group 467:  merge  transition  place  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	463 
    -- CP-element group 467: 	466 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	468 
    -- CP-element group 467:  members (2) 
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_919_PhiReqMerge
      -- CP-element group 467: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(467) <= OrReduce(convTranspose_CP_39_elements(463) & convTranspose_CP_39_elements(466));
    -- CP-element group 468:  fork  transition  place  input  output  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	467 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	222 
    -- CP-element group 468: 	223 
    -- CP-element group 468: 	225 
    -- CP-element group 468: 	227 
    -- CP-element group 468:  members (29) 
      -- CP-element group 468: 	 branch_block_stmt_32/merge_stmt_919__exit__
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950__entry__
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_update_start_
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resized_1
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scaled_1
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_computed_1
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/$exit
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/index_resize_req
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_resize_1/index_resize_ack
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/$exit
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/scale_rename_req
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_index_scale_1/scale_rename_ack
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_update_start
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Sample/req
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/array_obj_ref_932_final_index_sum_regn_Update/req
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/addr_of_933_complete/req
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_update_start_
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/$entry
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_934_to_assign_stmt_950/ptr_deref_936_Update/word_access_complete/word_0/cr
      -- CP-element group 468: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/$exit
      -- CP-element group 468: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/phi_stmt_920_ack
      -- 
    phi_stmt_920_ack_3537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_920_ack_0, ack => convTranspose_CP_39_elements(468)); -- 
    req_1763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(468), ack => array_obj_ref_932_index_offset_req_0); -- 
    req_1768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(468), ack => array_obj_ref_932_index_offset_req_1); -- 
    req_1783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(468), ack => addr_of_933_final_reg_req_1); -- 
    cr_1833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(468), ack => ptr_deref_936_store_0_req_1); -- 
    -- CP-element group 469:  merge  fork  transition  place  output  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	219 
    -- CP-element group 469: 	229 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	365 
    -- CP-element group 469: 	367 
    -- CP-element group 469: 	369 
    -- CP-element group 469: 	371 
    -- CP-element group 469: 	349 
    -- CP-element group 469: 	350 
    -- CP-element group 469: 	354 
    -- CP-element group 469: 	355 
    -- CP-element group 469: 	231 
    -- CP-element group 469: 	232 
    -- CP-element group 469: 	234 
    -- CP-element group 469: 	235 
    -- CP-element group 469: 	263 
    -- CP-element group 469: 	281 
    -- CP-element group 469: 	282 
    -- CP-element group 469: 	286 
    -- CP-element group 469: 	287 
    -- CP-element group 469: 	297 
    -- CP-element group 469: 	315 
    -- CP-element group 469: 	316 
    -- CP-element group 469: 	320 
    -- CP-element group 469: 	321 
    -- CP-element group 469: 	331 
    -- CP-element group 469:  members (76) 
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_update_start_
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_959__exit__
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192__entry__
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_Sample/req
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1048_Update/cr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block1_start_1013_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Sample/req
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Update/cr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block2_start_1069_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_update_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1055_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_update_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Sample/crr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/call_stmt_962_Update/ccr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_update_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_967_Update/cr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block0_start_969_Sample/req
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_update_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1104_Update/cr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_update_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1111_Update/cr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/WPIPE_Block3_start_1125_Sample/req
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_update_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1160_Update/cr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_update_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/type_cast_1167_Update/cr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block0_done_1182_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block1_done_1185_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block2_done_1188_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Sample/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/call_stmt_962_to_assign_stmt_1192/RPIPE_Block3_done_1191_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_959_PhiReqMerge
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_959_PhiAck/$entry
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_959_PhiAck/$exit
      -- CP-element group 469: 	 branch_block_stmt_32/merge_stmt_959_PhiAck/dummy
      -- 
    rr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1048_inst_req_0); -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => WPIPE_Block1_start_1013_inst_req_0); -- 
    cr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1048_inst_req_1); -- 
    req_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => WPIPE_Block2_start_1069_inst_req_0); -- 
    cr_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1055_inst_req_1); -- 
    rr_2242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1055_inst_req_0); -- 
    crr_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => call_stmt_962_call_req_0); -- 
    ccr_1869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => call_stmt_962_call_req_1); -- 
    cr_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_967_inst_req_1); -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => WPIPE_Block0_start_969_inst_req_0); -- 
    rr_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1104_inst_req_0); -- 
    cr_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1104_inst_req_1); -- 
    rr_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1111_inst_req_0); -- 
    cr_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1111_inst_req_1); -- 
    req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => WPIPE_Block3_start_1125_inst_req_0); -- 
    rr_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1160_inst_req_0); -- 
    cr_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1160_inst_req_1); -- 
    rr_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1167_inst_req_0); -- 
    cr_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => type_cast_1167_inst_req_1); -- 
    rr_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => RPIPE_Block0_done_1182_inst_req_0); -- 
    rr_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => RPIPE_Block1_done_1185_inst_req_0); -- 
    rr_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => RPIPE_Block2_done_1188_inst_req_0); -- 
    rr_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(469), ack => RPIPE_Block3_done_1191_inst_req_0); -- 
    convTranspose_CP_39_elements(469) <= OrReduce(convTranspose_CP_39_elements(219) & convTranspose_CP_39_elements(229));
    -- CP-element group 470:  transition  output  delay-element  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	400 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	474 
    -- CP-element group 470:  members (5) 
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph_forx_xbody419_PhiReq/$exit
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph_forx_xbody419_PhiReq/phi_stmt_1297/$exit
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/$exit
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1301_konst_delay_trans
      -- CP-element group 470: 	 branch_block_stmt_32/bbx_xnph_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_req
      -- 
    phi_stmt_1297_req_3583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1297_req_3583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(470), ack => phi_stmt_1297_req_0); -- 
    -- Element group convTranspose_CP_39_elements(470) is a control-delay.
    cp_element_470_delay: control_delay_element  generic map(name => " 470_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(400), ack => convTranspose_CP_39_elements(470), clk => clk, reset =>reset);
    -- CP-element group 471:  transition  input  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	448 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	473 
    -- CP-element group 471:  members (2) 
      -- CP-element group 471: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Sample/$exit
      -- CP-element group 471: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Sample/ra
      -- 
    ra_3603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1303_inst_ack_0, ack => convTranspose_CP_39_elements(471)); -- 
    -- CP-element group 472:  transition  input  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	448 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	473 
    -- CP-element group 472:  members (2) 
      -- CP-element group 472: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Update/$exit
      -- CP-element group 472: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/Update/ca
      -- 
    ca_3608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1303_inst_ack_1, ack => convTranspose_CP_39_elements(472)); -- 
    -- CP-element group 473:  join  transition  output  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	471 
    -- CP-element group 473: 	472 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473:  members (6) 
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_sources/type_cast_1303/SplitProtocol/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/forx_xbody419_forx_xbody419_PhiReq/phi_stmt_1297/phi_stmt_1297_req
      -- 
    phi_stmt_1297_req_3609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1297_req_3609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(473), ack => phi_stmt_1297_req_1); -- 
    convTranspose_cp_element_group_473: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_473"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(471) & convTranspose_CP_39_elements(472);
      gj_convTranspose_cp_element_group_473 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(473), clk => clk, reset => reset); --
    end block;
    -- CP-element group 474:  merge  transition  place  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	470 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474:  members (2) 
      -- CP-element group 474: 	 branch_block_stmt_32/merge_stmt_1296_PhiReqMerge
      -- CP-element group 474: 	 branch_block_stmt_32/merge_stmt_1296_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(474) <= OrReduce(convTranspose_CP_39_elements(470) & convTranspose_CP_39_elements(473));
    -- CP-element group 475:  fork  transition  place  input  output  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	474 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	401 
    -- CP-element group 475: 	402 
    -- CP-element group 475: 	404 
    -- CP-element group 475: 	406 
    -- CP-element group 475: 	408 
    -- CP-element group 475: 	410 
    -- CP-element group 475: 	412 
    -- CP-element group 475: 	414 
    -- CP-element group 475: 	416 
    -- CP-element group 475: 	418 
    -- CP-element group 475: 	420 
    -- CP-element group 475: 	422 
    -- CP-element group 475:  members (53) 
      -- CP-element group 475: 	 branch_block_stmt_32/merge_stmt_1296__exit__
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424__entry__
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_complete/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1328_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_complete/req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_final_index_sum_regn_Update/req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_final_index_sum_regn_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1368_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_final_index_sum_regn_Sample/req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1318_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_final_index_sum_regn_Sample/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_final_index_sum_regn_update_start
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_scale_1/scale_rename_ack
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1358_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_scale_1/scale_rename_req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/word_access_complete/word_0/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_scale_1/$exit
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/word_access_complete/word_0/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_scale_1/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1388_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/word_access_complete/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_resize_1/index_resize_ack
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_resize_1/index_resize_req
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/ptr_deref_1314_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_resize_1/$exit
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_resize_1/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_computed_1
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_scaled_1
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1348_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/array_obj_ref_1309_index_resized_1
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1378_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/addr_of_1310_update_start_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1311_to_assign_stmt_1424/type_cast_1338_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_32/merge_stmt_1296_PhiAck/$exit
      -- CP-element group 475: 	 branch_block_stmt_32/merge_stmt_1296_PhiAck/phi_stmt_1297_ack
      -- 
    phi_stmt_1297_ack_3614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1297_ack_0, ack => convTranspose_CP_39_elements(475)); -- 
    cr_3113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_1328_inst_req_1); -- 
    req_3035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => addr_of_1310_final_reg_req_1); -- 
    cr_3099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_1318_inst_req_1); -- 
    req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => array_obj_ref_1309_index_offset_req_1); -- 
    cr_3169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_1368_inst_req_1); -- 
    req_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => array_obj_ref_1309_index_offset_req_0); -- 
    cr_3197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_1388_inst_req_1); -- 
    cr_3155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_1358_inst_req_1); -- 
    cr_3080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => ptr_deref_1314_load_0_req_1); -- 
    cr_3141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_1348_inst_req_1); -- 
    cr_3183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_1378_inst_req_1); -- 
    cr_3127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(475), ack => type_cast_1338_inst_req_1); -- 
    -- CP-element group 476:  merge  transition  place  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	398 
    -- CP-element group 476: 	447 
    -- CP-element group 476: successors 
    -- CP-element group 476:  members (16) 
      -- CP-element group 476: 	 $exit
      -- CP-element group 476: 	 branch_block_stmt_32/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/branch_block_stmt_32__exit__
      -- CP-element group 476: 	 branch_block_stmt_32/merge_stmt_1433__exit__
      -- CP-element group 476: 	 branch_block_stmt_32/return__
      -- CP-element group 476: 	 branch_block_stmt_32/merge_stmt_1435__exit__
      -- CP-element group 476: 	 branch_block_stmt_32/merge_stmt_1433_PhiReqMerge
      -- CP-element group 476: 	 branch_block_stmt_32/merge_stmt_1433_PhiAck/$entry
      -- CP-element group 476: 	 branch_block_stmt_32/merge_stmt_1433_PhiAck/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/merge_stmt_1433_PhiAck/dummy
      -- CP-element group 476: 	 branch_block_stmt_32/return___PhiReq/$entry
      -- CP-element group 476: 	 branch_block_stmt_32/return___PhiReq/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/merge_stmt_1435_PhiReqMerge
      -- CP-element group 476: 	 branch_block_stmt_32/merge_stmt_1435_PhiAck/$entry
      -- CP-element group 476: 	 branch_block_stmt_32/merge_stmt_1435_PhiAck/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/merge_stmt_1435_PhiAck/dummy
      -- 
    convTranspose_CP_39_elements(476) <= OrReduce(convTranspose_CP_39_elements(398) & convTranspose_CP_39_elements(447));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar517_931_resized : std_logic_vector(13 downto 0);
    signal R_indvar517_931_scaled : std_logic_vector(13 downto 0);
    signal R_indvar531_687_resized : std_logic_vector(10 downto 0);
    signal R_indvar531_687_scaled : std_logic_vector(10 downto 0);
    signal R_indvar547_480_resized : std_logic_vector(13 downto 0);
    signal R_indvar547_480_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1308_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1308_scaled : std_logic_vector(13 downto 0);
    signal add108_333 : std_logic_vector(15 downto 0);
    signal add117_358 : std_logic_vector(15 downto 0);
    signal add126_383 : std_logic_vector(15 downto 0);
    signal add12_82 : std_logic_vector(15 downto 0);
    signal add135_408 : std_logic_vector(15 downto 0);
    signal add150_508 : std_logic_vector(63 downto 0);
    signal add156_526 : std_logic_vector(63 downto 0);
    signal add162_544 : std_logic_vector(63 downto 0);
    signal add168_562 : std_logic_vector(63 downto 0);
    signal add174_580 : std_logic_vector(63 downto 0);
    signal add180_598 : std_logic_vector(63 downto 0);
    signal add186_616 : std_logic_vector(63 downto 0);
    signal add206_715 : std_logic_vector(63 downto 0);
    signal add212_733 : std_logic_vector(63 downto 0);
    signal add218_751 : std_logic_vector(63 downto 0);
    signal add21_107 : std_logic_vector(15 downto 0);
    signal add224_769 : std_logic_vector(63 downto 0);
    signal add230_787 : std_logic_vector(63 downto 0);
    signal add236_805 : std_logic_vector(63 downto 0);
    signal add242_823 : std_logic_vector(63 downto 0);
    signal add30_132 : std_logic_vector(15 downto 0);
    signal add39_157 : std_logic_vector(15 downto 0);
    signal add48_182 : std_logic_vector(15 downto 0);
    signal add57_207 : std_logic_vector(15 downto 0);
    signal add74_247 : std_logic_vector(31 downto 0);
    signal add79_252 : std_logic_vector(31 downto 0);
    signal add99_308 : std_logic_vector(15 downto 0);
    signal add_57 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1309_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1309_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_481_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_688_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_688_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_932_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_932_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_690 : std_logic_vector(31 downto 0);
    signal arrayidx269_934 : std_logic_vector(31 downto 0);
    signal arrayidx424_1311 : std_logic_vector(31 downto 0);
    signal arrayidx_483 : std_logic_vector(31 downto 0);
    signal call101_311 : std_logic_vector(7 downto 0);
    signal call106_324 : std_logic_vector(7 downto 0);
    signal call10_73 : std_logic_vector(7 downto 0);
    signal call110_336 : std_logic_vector(7 downto 0);
    signal call115_349 : std_logic_vector(7 downto 0);
    signal call119_361 : std_logic_vector(7 downto 0);
    signal call124_374 : std_logic_vector(7 downto 0);
    signal call128_386 : std_logic_vector(7 downto 0);
    signal call133_399 : std_logic_vector(7 downto 0);
    signal call143_486 : std_logic_vector(7 downto 0);
    signal call147_499 : std_logic_vector(7 downto 0);
    signal call14_85 : std_logic_vector(7 downto 0);
    signal call153_517 : std_logic_vector(7 downto 0);
    signal call159_535 : std_logic_vector(7 downto 0);
    signal call165_553 : std_logic_vector(7 downto 0);
    signal call171_571 : std_logic_vector(7 downto 0);
    signal call177_589 : std_logic_vector(7 downto 0);
    signal call183_607 : std_logic_vector(7 downto 0);
    signal call199_693 : std_logic_vector(7 downto 0);
    signal call19_98 : std_logic_vector(7 downto 0);
    signal call203_706 : std_logic_vector(7 downto 0);
    signal call209_724 : std_logic_vector(7 downto 0);
    signal call215_742 : std_logic_vector(7 downto 0);
    signal call221_760 : std_logic_vector(7 downto 0);
    signal call227_778 : std_logic_vector(7 downto 0);
    signal call233_796 : std_logic_vector(7 downto 0);
    signal call239_814 : std_logic_vector(7 downto 0);
    signal call23_110 : std_logic_vector(7 downto 0);
    signal call275_962 : std_logic_vector(63 downto 0);
    signal call28_123 : std_logic_vector(7 downto 0);
    signal call2_48 : std_logic_vector(7 downto 0);
    signal call32_135 : std_logic_vector(7 downto 0);
    signal call346_1183 : std_logic_vector(15 downto 0);
    signal call348_1186 : std_logic_vector(15 downto 0);
    signal call350_1189 : std_logic_vector(15 downto 0);
    signal call352_1192 : std_logic_vector(15 downto 0);
    signal call354_1195 : std_logic_vector(63 downto 0);
    signal call37_148 : std_logic_vector(7 downto 0);
    signal call41_160 : std_logic_vector(7 downto 0);
    signal call46_173 : std_logic_vector(7 downto 0);
    signal call50_185 : std_logic_vector(7 downto 0);
    signal call55_198 : std_logic_vector(7 downto 0);
    signal call5_60 : std_logic_vector(7 downto 0);
    signal call92_286 : std_logic_vector(7 downto 0);
    signal call97_299 : std_logic_vector(7 downto 0);
    signal call_35 : std_logic_vector(7 downto 0);
    signal cmp194501_430 : std_logic_vector(0 downto 0);
    signal cmp264497_875 : std_logic_vector(0 downto 0);
    signal cmp505_415 : std_logic_vector(0 downto 0);
    signal conv104_315 : std_logic_vector(15 downto 0);
    signal conv107_328 : std_logic_vector(15 downto 0);
    signal conv113_340 : std_logic_vector(15 downto 0);
    signal conv116_353 : std_logic_vector(15 downto 0);
    signal conv11_77 : std_logic_vector(15 downto 0);
    signal conv122_365 : std_logic_vector(15 downto 0);
    signal conv125_378 : std_logic_vector(15 downto 0);
    signal conv131_390 : std_logic_vector(15 downto 0);
    signal conv134_403 : std_logic_vector(15 downto 0);
    signal conv144_490 : std_logic_vector(63 downto 0);
    signal conv149_503 : std_logic_vector(63 downto 0);
    signal conv155_521 : std_logic_vector(63 downto 0);
    signal conv161_539 : std_logic_vector(63 downto 0);
    signal conv167_557 : std_logic_vector(63 downto 0);
    signal conv173_575 : std_logic_vector(63 downto 0);
    signal conv179_593 : std_logic_vector(63 downto 0);
    signal conv17_89 : std_logic_vector(15 downto 0);
    signal conv185_611 : std_logic_vector(63 downto 0);
    signal conv1_39 : std_logic_vector(15 downto 0);
    signal conv200_697 : std_logic_vector(63 downto 0);
    signal conv205_710 : std_logic_vector(63 downto 0);
    signal conv20_102 : std_logic_vector(15 downto 0);
    signal conv211_728 : std_logic_vector(63 downto 0);
    signal conv217_746 : std_logic_vector(63 downto 0);
    signal conv223_764 : std_logic_vector(63 downto 0);
    signal conv229_782 : std_logic_vector(63 downto 0);
    signal conv235_800 : std_logic_vector(63 downto 0);
    signal conv241_818 : std_logic_vector(63 downto 0);
    signal conv253_851 : std_logic_vector(31 downto 0);
    signal conv255_855 : std_logic_vector(31 downto 0);
    signal conv258_859 : std_logic_vector(31 downto 0);
    signal conv26_114 : std_logic_vector(15 downto 0);
    signal conv276_968 : std_logic_vector(63 downto 0);
    signal conv29_127 : std_logic_vector(15 downto 0);
    signal conv305_1049 : std_logic_vector(15 downto 0);
    signal conv307_1056 : std_logic_vector(15 downto 0);
    signal conv322_1105 : std_logic_vector(15 downto 0);
    signal conv324_1112 : std_logic_vector(15 downto 0);
    signal conv339_1161 : std_logic_vector(15 downto 0);
    signal conv341_1168 : std_logic_vector(15 downto 0);
    signal conv355_1200 : std_logic_vector(63 downto 0);
    signal conv35_139 : std_logic_vector(15 downto 0);
    signal conv361_1209 : std_logic_vector(7 downto 0);
    signal conv367_1219 : std_logic_vector(7 downto 0);
    signal conv373_1229 : std_logic_vector(7 downto 0);
    signal conv379_1239 : std_logic_vector(7 downto 0);
    signal conv38_152 : std_logic_vector(15 downto 0);
    signal conv3_52 : std_logic_vector(15 downto 0);
    signal conv429_1319 : std_logic_vector(7 downto 0);
    signal conv435_1329 : std_logic_vector(7 downto 0);
    signal conv441_1339 : std_logic_vector(7 downto 0);
    signal conv447_1349 : std_logic_vector(7 downto 0);
    signal conv44_164 : std_logic_vector(15 downto 0);
    signal conv453_1359 : std_logic_vector(7 downto 0);
    signal conv459_1369 : std_logic_vector(7 downto 0);
    signal conv465_1379 : std_logic_vector(7 downto 0);
    signal conv471_1389 : std_logic_vector(7 downto 0);
    signal conv47_177 : std_logic_vector(15 downto 0);
    signal conv53_189 : std_logic_vector(15 downto 0);
    signal conv56_202 : std_logic_vector(15 downto 0);
    signal conv61_211 : std_logic_vector(31 downto 0);
    signal conv63_215 : std_logic_vector(31 downto 0);
    signal conv65_219 : std_logic_vector(31 downto 0);
    signal conv82_256 : std_logic_vector(31 downto 0);
    signal conv84_260 : std_logic_vector(31 downto 0);
    signal conv87_264 : std_logic_vector(31 downto 0);
    signal conv8_64 : std_logic_vector(15 downto 0);
    signal conv90_268 : std_logic_vector(31 downto 0);
    signal conv95_290 : std_logic_vector(15 downto 0);
    signal conv98_303 : std_logic_vector(15 downto 0);
    signal exitcond1_1424 : std_logic_vector(0 downto 0);
    signal exitcond2_838 : std_logic_vector(0 downto 0);
    signal exitcond3_631 : std_logic_vector(0 downto 0);
    signal exitcond_950 : std_logic_vector(0 downto 0);
    signal iNsTr_14_241 : std_logic_vector(31 downto 0);
    signal iNsTr_186_1281 : std_logic_vector(63 downto 0);
    signal iNsTr_26_453 : std_logic_vector(63 downto 0);
    signal iNsTr_39_660 : std_logic_vector(63 downto 0);
    signal iNsTr_53_904 : std_logic_vector(63 downto 0);
    signal indvar517_920 : std_logic_vector(63 downto 0);
    signal indvar531_676 : std_logic_vector(63 downto 0);
    signal indvar547_469 : std_logic_vector(63 downto 0);
    signal indvar_1297 : std_logic_vector(63 downto 0);
    signal indvarx_xnext518_945 : std_logic_vector(63 downto 0);
    signal indvarx_xnext532_833 : std_logic_vector(63 downto 0);
    signal indvarx_xnext548_626 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1419 : std_logic_vector(63 downto 0);
    signal mul256_864 : std_logic_vector(31 downto 0);
    signal mul259_869 : std_logic_vector(31 downto 0);
    signal mul66_229 : std_logic_vector(31 downto 0);
    signal mul85_273 : std_logic_vector(31 downto 0);
    signal mul88_278 : std_logic_vector(31 downto 0);
    signal mul91_283 : std_logic_vector(31 downto 0);
    signal mul_224 : std_logic_vector(31 downto 0);
    signal ptr_deref_1314_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1314_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1314_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1314_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1314_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_618_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_618_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_618_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_618_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_618_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_618_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_825_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_825_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_825_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_825_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_825_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_825_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_936_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_936_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_936_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_936_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_936_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_936_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_321 : std_logic_vector(15 downto 0);
    signal shl114_346 : std_logic_vector(15 downto 0);
    signal shl123_371 : std_logic_vector(15 downto 0);
    signal shl132_396 : std_logic_vector(15 downto 0);
    signal shl146_496 : std_logic_vector(63 downto 0);
    signal shl152_514 : std_logic_vector(63 downto 0);
    signal shl158_532 : std_logic_vector(63 downto 0);
    signal shl164_550 : std_logic_vector(63 downto 0);
    signal shl170_568 : std_logic_vector(63 downto 0);
    signal shl176_586 : std_logic_vector(63 downto 0);
    signal shl182_604 : std_logic_vector(63 downto 0);
    signal shl18_95 : std_logic_vector(15 downto 0);
    signal shl202_703 : std_logic_vector(63 downto 0);
    signal shl208_721 : std_logic_vector(63 downto 0);
    signal shl214_739 : std_logic_vector(63 downto 0);
    signal shl220_757 : std_logic_vector(63 downto 0);
    signal shl226_775 : std_logic_vector(63 downto 0);
    signal shl232_793 : std_logic_vector(63 downto 0);
    signal shl238_811 : std_logic_vector(63 downto 0);
    signal shl27_120 : std_logic_vector(15 downto 0);
    signal shl36_145 : std_logic_vector(15 downto 0);
    signal shl45_170 : std_logic_vector(15 downto 0);
    signal shl54_195 : std_logic_vector(15 downto 0);
    signal shl96_296 : std_logic_vector(15 downto 0);
    signal shl9_70 : std_logic_vector(15 downto 0);
    signal shl_45 : std_logic_vector(15 downto 0);
    signal shr304_1045 : std_logic_vector(31 downto 0);
    signal shr321_1101 : std_logic_vector(31 downto 0);
    signal shr338_1157 : std_logic_vector(31 downto 0);
    signal shr364_1215 : std_logic_vector(63 downto 0);
    signal shr370_1225 : std_logic_vector(63 downto 0);
    signal shr376_1235 : std_logic_vector(63 downto 0);
    signal shr432_1325 : std_logic_vector(63 downto 0);
    signal shr438_1335 : std_logic_vector(63 downto 0);
    signal shr444_1345 : std_logic_vector(63 downto 0);
    signal shr450_1355 : std_logic_vector(63 downto 0);
    signal shr456_1365 : std_logic_vector(63 downto 0);
    signal shr462_1375 : std_logic_vector(63 downto 0);
    signal shr468_1385 : std_logic_vector(63 downto 0);
    signal shr_235 : std_logic_vector(31 downto 0);
    signal sub_1205 : std_logic_vector(63 downto 0);
    signal tmp425_1315 : std_logic_vector(63 downto 0);
    signal tmp512_1265 : std_logic_vector(31 downto 0);
    signal tmp512x_xop_1277 : std_logic_vector(31 downto 0);
    signal tmp513_1271 : std_logic_vector(0 downto 0);
    signal tmp516_1294 : std_logic_vector(63 downto 0);
    signal tmp524_888 : std_logic_vector(31 downto 0);
    signal tmp524x_xop_900 : std_logic_vector(31 downto 0);
    signal tmp525_894 : std_logic_vector(0 downto 0);
    signal tmp529_917 : std_logic_vector(63 downto 0);
    signal tmp540_644 : std_logic_vector(31 downto 0);
    signal tmp540x_xop_656 : std_logic_vector(31 downto 0);
    signal tmp541_650 : std_logic_vector(0 downto 0);
    signal tmp545_673 : std_logic_vector(63 downto 0);
    signal tmp554x_xop_449 : std_logic_vector(31 downto 0);
    signal tmp555_443 : std_logic_vector(0 downto 0);
    signal tmp559_466 : std_logic_vector(63 downto 0);
    signal type_cast_1002_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1043_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1099_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1155_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_118_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1198_wire : std_logic_vector(63 downto 0);
    signal type_cast_1213_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1223_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1233_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1263_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1269_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1275_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1285_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1292_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1301_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1303_wire : std_logic_vector(63 downto 0);
    signal type_cast_1323_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1333_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1343_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1353_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1363_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1373_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1383_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1417_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_143_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_168_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_193_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_233_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_239_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_245_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_294_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_319_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_344_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_369_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_394_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_412_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_428_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_43_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_441_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_447_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_464_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_473_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_475_wire : std_logic_vector(63 downto 0);
    signal type_cast_494_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_530_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_548_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_584_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_602_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_624_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_642_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_648_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_664_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_671_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_679_wire : std_logic_vector(63 downto 0);
    signal type_cast_682_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_68_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_701_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_719_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_737_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_773_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_791_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_809_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_831_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_873_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_886_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_892_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_898_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_908_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_915_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_923_wire : std_logic_vector(63 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_938_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_93_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_943_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_966_wire : std_logic_vector(63 downto 0);
    signal type_cast_998_wire_constant : std_logic_vector(15 downto 0);
    signal xx_xop561_910 : std_logic_vector(63 downto 0);
    signal xx_xop562_666 : std_logic_vector(63 downto 0);
    signal xx_xop563_459 : std_logic_vector(63 downto 0);
    signal xx_xop_1287 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1309_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1309_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1309_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1309_resized_base_address <= "00000000000000";
    array_obj_ref_481_constant_part_of_offset <= "00000000000000";
    array_obj_ref_481_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_481_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_481_resized_base_address <= "00000000000000";
    array_obj_ref_688_constant_part_of_offset <= "00000100010";
    array_obj_ref_688_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_688_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_688_resized_base_address <= "00000000000";
    array_obj_ref_932_constant_part_of_offset <= "00000000000000";
    array_obj_ref_932_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_932_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_932_resized_base_address <= "00000000000000";
    ptr_deref_1314_word_offset_0 <= "00000000000000";
    ptr_deref_618_word_offset_0 <= "00000000000000";
    ptr_deref_825_word_offset_0 <= "00000000000";
    ptr_deref_936_word_offset_0 <= "00000000000000";
    type_cast_1002_wire_constant <= "0000000000000000";
    type_cast_1043_wire_constant <= "00000000000000000000000000010010";
    type_cast_1099_wire_constant <= "00000000000000000000000000010001";
    type_cast_1155_wire_constant <= "00000000000000000000000000010000";
    type_cast_118_wire_constant <= "0000000000001000";
    type_cast_1213_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1223_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1233_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1263_wire_constant <= "00000000000000000000000000000010";
    type_cast_1269_wire_constant <= "00000000000000000000000000000001";
    type_cast_1275_wire_constant <= "11111111111111111111111111111111";
    type_cast_1285_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1292_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1301_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1323_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1333_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1343_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1353_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1363_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1373_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1383_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1417_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_143_wire_constant <= "0000000000001000";
    type_cast_168_wire_constant <= "0000000000001000";
    type_cast_193_wire_constant <= "0000000000001000";
    type_cast_233_wire_constant <= "00000000000000000000000000000010";
    type_cast_239_wire_constant <= "00000000000000000000000000000001";
    type_cast_245_wire_constant <= "01111111111111111111111111111110";
    type_cast_294_wire_constant <= "0000000000001000";
    type_cast_319_wire_constant <= "0000000000001000";
    type_cast_344_wire_constant <= "0000000000001000";
    type_cast_369_wire_constant <= "0000000000001000";
    type_cast_394_wire_constant <= "0000000000001000";
    type_cast_412_wire_constant <= "00000000000000000000000000000011";
    type_cast_428_wire_constant <= "00000000000000000000000000000011";
    type_cast_43_wire_constant <= "0000000000001000";
    type_cast_441_wire_constant <= "00000000000000000000000000000001";
    type_cast_447_wire_constant <= "11111111111111111111111111111111";
    type_cast_457_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_464_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_473_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_494_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_512_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_530_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_548_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_566_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_584_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_602_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_624_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_642_wire_constant <= "00000000000000000000000000000010";
    type_cast_648_wire_constant <= "00000000000000000000000000000001";
    type_cast_654_wire_constant <= "11111111111111111111111111111111";
    type_cast_664_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_671_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_682_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_68_wire_constant <= "0000000000001000";
    type_cast_701_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_719_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_737_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_755_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_773_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_791_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_809_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_831_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_873_wire_constant <= "00000000000000000000000000000011";
    type_cast_886_wire_constant <= "00000000000000000000000000000010";
    type_cast_892_wire_constant <= "00000000000000000000000000000001";
    type_cast_898_wire_constant <= "11111111111111111111111111111111";
    type_cast_908_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_915_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_926_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_938_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_93_wire_constant <= "0000000000001000";
    type_cast_943_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_998_wire_constant <= "0000000000000000";
    phi_stmt_1297: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1301_wire_constant & type_cast_1303_wire;
      req <= phi_stmt_1297_req_0 & phi_stmt_1297_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1297",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1297_ack_0,
          idata => idata,
          odata => indvar_1297,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1297
    phi_stmt_469: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_473_wire_constant & type_cast_475_wire;
      req <= phi_stmt_469_req_0 & phi_stmt_469_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_469",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_469_ack_0,
          idata => idata,
          odata => indvar547_469,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_469
    phi_stmt_676: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_679_wire & type_cast_682_wire_constant;
      req <= phi_stmt_676_req_0 & phi_stmt_676_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_676",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_676_ack_0,
          idata => idata,
          odata => indvar531_676,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_676
    phi_stmt_920: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_923_wire & type_cast_926_wire_constant;
      req <= phi_stmt_920_req_0 & phi_stmt_920_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_920",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_920_ack_0,
          idata => idata,
          odata => indvar517_920,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_920
    -- flow-through select operator MUX_1293_inst
    tmp516_1294 <= xx_xop_1287 when (tmp513_1271(0) /=  '0') else type_cast_1292_wire_constant;
    -- flow-through select operator MUX_465_inst
    tmp559_466 <= xx_xop563_459 when (tmp555_443(0) /=  '0') else type_cast_464_wire_constant;
    -- flow-through select operator MUX_672_inst
    tmp545_673 <= xx_xop562_666 when (tmp541_650(0) /=  '0') else type_cast_671_wire_constant;
    -- flow-through select operator MUX_916_inst
    tmp529_917 <= xx_xop561_910 when (tmp525_894(0) /=  '0') else type_cast_915_wire_constant;
    addr_of_1310_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1310_final_reg_req_0;
      addr_of_1310_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1310_final_reg_req_1;
      addr_of_1310_final_reg_ack_1<= rack(0);
      addr_of_1310_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1310_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1309_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx424_1311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_482_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_482_final_reg_req_0;
      addr_of_482_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_482_final_reg_req_1;
      addr_of_482_final_reg_ack_1<= rack(0);
      addr_of_482_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_482_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_481_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_689_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_689_final_reg_req_0;
      addr_of_689_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_689_final_reg_req_1;
      addr_of_689_final_reg_ack_1<= rack(0);
      addr_of_689_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_689_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_688_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_933_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_933_final_reg_req_0;
      addr_of_933_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_933_final_reg_req_1;
      addr_of_933_final_reg_ack_1<= rack(0);
      addr_of_933_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_933_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_932_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_934,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_101_inst_req_0;
      type_cast_101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_101_inst_req_1;
      type_cast_101_inst_ack_1<= rack(0);
      type_cast_101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_98,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1048_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1048_inst_req_0;
      type_cast_1048_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1048_inst_req_1;
      type_cast_1048_inst_ack_1<= rack(0);
      type_cast_1048_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1048_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr304_1045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1049,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1055_inst_req_0;
      type_cast_1055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1055_inst_req_1;
      type_cast_1055_inst_ack_1<= rack(0);
      type_cast_1055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1055_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv307_1056,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1104_inst_req_0;
      type_cast_1104_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1104_inst_req_1;
      type_cast_1104_inst_ack_1<= rack(0);
      type_cast_1104_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1104_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr321_1101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1105,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1111_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1111_inst_req_0;
      type_cast_1111_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1111_inst_req_1;
      type_cast_1111_inst_ack_1<= rack(0);
      type_cast_1111_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1111_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add74_247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv324_1112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_113_inst_req_0;
      type_cast_113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_113_inst_req_1;
      type_cast_113_inst_ack_1<= rack(0);
      type_cast_113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_110,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1160_inst_req_0;
      type_cast_1160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1160_inst_req_1;
      type_cast_1160_inst_ack_1<= rack(0);
      type_cast_1160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv339_1161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1167_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1167_inst_req_0;
      type_cast_1167_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1167_inst_req_1;
      type_cast_1167_inst_ack_1<= rack(0);
      type_cast_1167_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1167_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79_252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1199_inst_req_0;
      type_cast_1199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1199_inst_req_1;
      type_cast_1199_inst_ack_1<= rack(0);
      type_cast_1199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1198_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv355_1200,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1208_inst_req_0;
      type_cast_1208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1208_inst_req_1;
      type_cast_1208_inst_ack_1<= rack(0);
      type_cast_1208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1205,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv361_1209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1218_inst_req_0;
      type_cast_1218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1218_inst_req_1;
      type_cast_1218_inst_ack_1<= rack(0);
      type_cast_1218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr364_1215,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv367_1219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1228_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1228_inst_req_0;
      type_cast_1228_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1228_inst_req_1;
      type_cast_1228_inst_ack_1<= rack(0);
      type_cast_1228_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1228_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr370_1225,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv373_1229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr376_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv379_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_126_inst_req_0;
      type_cast_126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_126_inst_req_1;
      type_cast_126_inst_ack_1<= rack(0);
      type_cast_126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1280_inst_req_0;
      type_cast_1280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1280_inst_req_1;
      type_cast_1280_inst_ack_1<= rack(0);
      type_cast_1280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1280_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp512x_xop_1277,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_186_1281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1303_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1303_inst_req_0;
      type_cast_1303_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1303_inst_req_1;
      type_cast_1303_inst_ack_1<= rack(0);
      type_cast_1303_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1303_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1303_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1318_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1318_inst_req_0;
      type_cast_1318_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1318_inst_req_1;
      type_cast_1318_inst_ack_1<= rack(0);
      type_cast_1318_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1318_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp425_1315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv429_1319,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1328_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1328_inst_req_0;
      type_cast_1328_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1328_inst_req_1;
      type_cast_1328_inst_ack_1<= rack(0);
      type_cast_1328_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1328_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr432_1325,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv435_1329,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1338_inst_req_0;
      type_cast_1338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1338_inst_req_1;
      type_cast_1338_inst_ack_1<= rack(0);
      type_cast_1338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr438_1335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv441_1339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1348_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1348_inst_req_0;
      type_cast_1348_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1348_inst_req_1;
      type_cast_1348_inst_ack_1<= rack(0);
      type_cast_1348_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1348_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr444_1345,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv447_1349,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1358_inst_req_0;
      type_cast_1358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1358_inst_req_1;
      type_cast_1358_inst_ack_1<= rack(0);
      type_cast_1358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr450_1355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv453_1359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1368_inst_req_0;
      type_cast_1368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1368_inst_req_1;
      type_cast_1368_inst_ack_1<= rack(0);
      type_cast_1368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr456_1365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv459_1369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1378_inst_req_0;
      type_cast_1378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1378_inst_req_1;
      type_cast_1378_inst_ack_1<= rack(0);
      type_cast_1378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr462_1375,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv465_1379,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1388_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1388_inst_req_0;
      type_cast_1388_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1388_inst_req_1;
      type_cast_1388_inst_ack_1<= rack(0);
      type_cast_1388_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1388_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr468_1385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv471_1389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_138_inst_req_0;
      type_cast_138_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_138_inst_req_1;
      type_cast_138_inst_ack_1<= rack(0);
      type_cast_138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_151_inst_req_0;
      type_cast_151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_151_inst_req_1;
      type_cast_151_inst_ack_1<= rack(0);
      type_cast_151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_152,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_163_inst_req_0;
      type_cast_163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_163_inst_req_1;
      type_cast_163_inst_ack_1<= rack(0);
      type_cast_163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_176_inst_req_0;
      type_cast_176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_176_inst_req_1;
      type_cast_176_inst_ack_1<= rack(0);
      type_cast_176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_188_inst_req_0;
      type_cast_188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_188_inst_req_1;
      type_cast_188_inst_ack_1<= rack(0);
      type_cast_188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_201_inst_req_0;
      type_cast_201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_201_inst_req_1;
      type_cast_201_inst_ack_1<= rack(0);
      type_cast_201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_210_inst_req_0;
      type_cast_210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_210_inst_req_1;
      type_cast_210_inst_ack_1<= rack(0);
      type_cast_210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_57,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_214_inst_req_0;
      type_cast_214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_214_inst_req_1;
      type_cast_214_inst_ack_1<= rack(0);
      type_cast_214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_82,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_218_inst_req_0;
      type_cast_218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_218_inst_req_1;
      type_cast_218_inst_ack_1<= rack(0);
      type_cast_218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_255_inst_req_0;
      type_cast_255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_255_inst_req_1;
      type_cast_255_inst_ack_1<= rack(0);
      type_cast_255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_259_inst_req_0;
      type_cast_259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_259_inst_req_1;
      type_cast_259_inst_ack_1<= rack(0);
      type_cast_259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_260,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_263_inst_req_0;
      type_cast_263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_263_inst_req_1;
      type_cast_263_inst_ack_1<= rack(0);
      type_cast_263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_182,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_264,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_267_inst_req_0;
      type_cast_267_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_267_inst_req_1;
      type_cast_267_inst_ack_1<= rack(0);
      type_cast_267_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_267_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_268,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_289_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_289_inst_req_0;
      type_cast_289_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_289_inst_req_1;
      type_cast_289_inst_ack_1<= rack(0);
      type_cast_289_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_289_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_290,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_302_inst_req_0;
      type_cast_302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_302_inst_req_1;
      type_cast_302_inst_ack_1<= rack(0);
      type_cast_302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_314_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_314_inst_req_0;
      type_cast_314_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_314_inst_req_1;
      type_cast_314_inst_ack_1<= rack(0);
      type_cast_314_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_314_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_315,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_327_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_327_inst_req_0;
      type_cast_327_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_327_inst_req_1;
      type_cast_327_inst_ack_1<= rack(0);
      type_cast_327_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_327_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_324,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_328,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_339_inst_req_0;
      type_cast_339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_339_inst_req_1;
      type_cast_339_inst_ack_1<= rack(0);
      type_cast_339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_352_inst_req_0;
      type_cast_352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_352_inst_req_1;
      type_cast_352_inst_ack_1<= rack(0);
      type_cast_352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_364_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_364_inst_req_0;
      type_cast_364_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_364_inst_req_1;
      type_cast_364_inst_ack_1<= rack(0);
      type_cast_364_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_364_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_361,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_365,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_377_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_377_inst_req_0;
      type_cast_377_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_377_inst_req_1;
      type_cast_377_inst_ack_1<= rack(0);
      type_cast_377_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_377_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_374,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_378,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_389_inst_req_0;
      type_cast_389_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_389_inst_req_1;
      type_cast_389_inst_ack_1<= rack(0);
      type_cast_389_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_390,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_38_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_38_inst_req_0;
      type_cast_38_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_38_inst_req_1;
      type_cast_38_inst_ack_1<= rack(0);
      type_cast_38_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_38_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_39,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_402_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_402_inst_req_0;
      type_cast_402_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_402_inst_req_1;
      type_cast_402_inst_ack_1<= rack(0);
      type_cast_402_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_402_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_399,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_452_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_452_inst_req_0;
      type_cast_452_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_452_inst_req_1;
      type_cast_452_inst_ack_1<= rack(0);
      type_cast_452_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_452_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp554x_xop_449,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_453,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_475_inst_req_0;
      type_cast_475_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_475_inst_req_1;
      type_cast_475_inst_ack_1<= rack(0);
      type_cast_475_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_475_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext548_626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_475_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_489_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_489_inst_req_0;
      type_cast_489_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_489_inst_req_1;
      type_cast_489_inst_ack_1<= rack(0);
      type_cast_489_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_489_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_486,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_490,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_502_inst_req_0;
      type_cast_502_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_502_inst_req_1;
      type_cast_502_inst_ack_1<= rack(0);
      type_cast_502_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_502_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_499,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_503,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_51_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_51_inst_req_0;
      type_cast_51_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_51_inst_req_1;
      type_cast_51_inst_ack_1<= rack(0);
      type_cast_51_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_51_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_48,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_52,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_520_inst_req_0;
      type_cast_520_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_520_inst_req_1;
      type_cast_520_inst_ack_1<= rack(0);
      type_cast_520_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_520_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_538_inst_req_0;
      type_cast_538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_538_inst_req_1;
      type_cast_538_inst_ack_1<= rack(0);
      type_cast_538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_556_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_556_inst_req_0;
      type_cast_556_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_556_inst_req_1;
      type_cast_556_inst_ack_1<= rack(0);
      type_cast_556_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_556_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_553,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_557,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_574_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_574_inst_req_0;
      type_cast_574_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_574_inst_req_1;
      type_cast_574_inst_ack_1<= rack(0);
      type_cast_574_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_574_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_571,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_575,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_592_inst_req_0;
      type_cast_592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_592_inst_req_1;
      type_cast_592_inst_ack_1<= rack(0);
      type_cast_592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_610_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_610_inst_req_0;
      type_cast_610_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_610_inst_req_1;
      type_cast_610_inst_ack_1<= rack(0);
      type_cast_610_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_610_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_611,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_63_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_63_inst_req_0;
      type_cast_63_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_63_inst_req_1;
      type_cast_63_inst_ack_1<= rack(0);
      type_cast_63_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_63_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_60,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_659_inst_req_0;
      type_cast_659_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_659_inst_req_1;
      type_cast_659_inst_ack_1<= rack(0);
      type_cast_659_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_659_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp540x_xop_656,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_660,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_679_inst_req_0;
      type_cast_679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_679_inst_req_1;
      type_cast_679_inst_ack_1<= rack(0);
      type_cast_679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_679_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext532_833,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_679_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_696_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_696_inst_req_0;
      type_cast_696_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_696_inst_req_1;
      type_cast_696_inst_ack_1<= rack(0);
      type_cast_696_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_696_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_693,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_697,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_709_inst_req_0;
      type_cast_709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_709_inst_req_1;
      type_cast_709_inst_ack_1<= rack(0);
      type_cast_709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_706,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_727_inst_req_0;
      type_cast_727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_727_inst_req_1;
      type_cast_727_inst_ack_1<= rack(0);
      type_cast_727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_724,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_745_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_745_inst_req_0;
      type_cast_745_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_745_inst_req_1;
      type_cast_745_inst_ack_1<= rack(0);
      type_cast_745_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_745_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_742,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_746,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_763_inst_req_0;
      type_cast_763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_763_inst_req_1;
      type_cast_763_inst_ack_1<= rack(0);
      type_cast_763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_760,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_73,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_781_inst_req_0;
      type_cast_781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_781_inst_req_1;
      type_cast_781_inst_ack_1<= rack(0);
      type_cast_781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_781_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_799_inst_req_0;
      type_cast_799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_799_inst_req_1;
      type_cast_799_inst_ack_1<= rack(0);
      type_cast_799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_800,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_817_inst_req_0;
      type_cast_817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_817_inst_req_1;
      type_cast_817_inst_ack_1<= rack(0);
      type_cast_817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_850_inst_req_0;
      type_cast_850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_850_inst_req_1;
      type_cast_850_inst_ack_1<= rack(0);
      type_cast_850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_851,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_854_inst_req_0;
      type_cast_854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_854_inst_req_1;
      type_cast_854_inst_ack_1<= rack(0);
      type_cast_854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_858_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_858_inst_req_0;
      type_cast_858_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_858_inst_req_1;
      type_cast_858_inst_ack_1<= rack(0);
      type_cast_858_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_858_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_408,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_859,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_88_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_88_inst_req_0;
      type_cast_88_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_88_inst_req_1;
      type_cast_88_inst_ack_1<= rack(0);
      type_cast_88_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_88_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_85,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_89,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_903_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_903_inst_req_0;
      type_cast_903_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_903_inst_req_1;
      type_cast_903_inst_ack_1<= rack(0);
      type_cast_903_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_903_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp524x_xop_900,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_904,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_923_inst_req_0;
      type_cast_923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_923_inst_req_1;
      type_cast_923_inst_ack_1<= rack(0);
      type_cast_923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext518_945,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_923_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_967_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_967_inst_req_0;
      type_cast_967_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_967_inst_req_1;
      type_cast_967_inst_ack_1<= rack(0);
      type_cast_967_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_967_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_966_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_968,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1309_index_1_rename
    process(R_indvar_1308_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1308_resized;
      ov(13 downto 0) := iv;
      R_indvar_1308_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1309_index_1_resize
    process(indvar_1297) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1297;
      ov := iv(13 downto 0);
      R_indvar_1308_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1309_root_address_inst
    process(array_obj_ref_1309_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1309_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1309_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_481_index_1_rename
    process(R_indvar547_480_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar547_480_resized;
      ov(13 downto 0) := iv;
      R_indvar547_480_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_481_index_1_resize
    process(indvar547_469) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar547_469;
      ov := iv(13 downto 0);
      R_indvar547_480_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_481_root_address_inst
    process(array_obj_ref_481_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_481_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_481_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_688_index_1_rename
    process(R_indvar531_687_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar531_687_resized;
      ov(10 downto 0) := iv;
      R_indvar531_687_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_688_index_1_resize
    process(indvar531_676) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar531_676;
      ov := iv(10 downto 0);
      R_indvar531_687_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_688_root_address_inst
    process(array_obj_ref_688_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_688_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_688_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_932_index_1_rename
    process(R_indvar517_931_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar517_931_resized;
      ov(13 downto 0) := iv;
      R_indvar517_931_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_932_index_1_resize
    process(indvar517_920) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar517_920;
      ov := iv(13 downto 0);
      R_indvar517_931_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_932_root_address_inst
    process(array_obj_ref_932_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_932_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_932_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1314_addr_0
    process(ptr_deref_1314_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1314_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1314_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1314_base_resize
    process(arrayidx424_1311) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx424_1311;
      ov := iv(13 downto 0);
      ptr_deref_1314_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1314_gather_scatter
    process(ptr_deref_1314_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1314_data_0;
      ov(63 downto 0) := iv;
      tmp425_1315 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1314_root_address_inst
    process(ptr_deref_1314_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1314_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1314_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_addr_0
    process(ptr_deref_618_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_618_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_618_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_base_resize
    process(arrayidx_483) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_483;
      ov := iv(13 downto 0);
      ptr_deref_618_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_gather_scatter
    process(add186_616) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_616;
      ov(63 downto 0) := iv;
      ptr_deref_618_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_618_root_address_inst
    process(ptr_deref_618_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_618_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_618_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_addr_0
    process(ptr_deref_825_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_825_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_825_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_base_resize
    process(arrayidx246_690) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_690;
      ov := iv(10 downto 0);
      ptr_deref_825_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_gather_scatter
    process(add242_823) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_823;
      ov(63 downto 0) := iv;
      ptr_deref_825_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_825_root_address_inst
    process(ptr_deref_825_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_825_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_825_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_addr_0
    process(ptr_deref_936_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_936_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_936_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_base_resize
    process(arrayidx269_934) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_934;
      ov := iv(13 downto 0);
      ptr_deref_936_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_gather_scatter
    process(type_cast_938_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_938_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_936_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_root_address_inst
    process(ptr_deref_936_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_936_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_936_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1253_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264497_875;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1253_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1253_branch_req_0,
          ack0 => if_stmt_1253_branch_ack_0,
          ack1 => if_stmt_1253_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1425_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1424;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1425_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1425_branch_req_0,
          ack0 => if_stmt_1425_branch_ack_0,
          ack1 => if_stmt_1425_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_416_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp505_415;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_416_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_416_branch_req_0,
          ack0 => if_stmt_416_branch_ack_0,
          ack1 => if_stmt_416_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_431_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194501_430;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_431_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_431_branch_req_0,
          ack0 => if_stmt_431_branch_ack_0,
          ack1 => if_stmt_431_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_632_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_631;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_632_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_632_branch_req_0,
          ack0 => if_stmt_632_branch_ack_0,
          ack1 => if_stmt_632_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_839_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_838;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_839_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_839_branch_req_0,
          ack0 => if_stmt_839_branch_ack_0,
          ack1 => if_stmt_839_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_876_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264497_875;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_876_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_876_branch_req_0,
          ack0 => if_stmt_876_branch_ack_0,
          ack1 => if_stmt_876_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_951_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_950;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_951_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_951_branch_req_0,
          ack0 => if_stmt_951_branch_ack_0,
          ack1 => if_stmt_951_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1276_inst
    process(tmp512_1265) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp512_1265, type_cast_1275_wire_constant, tmp_var);
      tmp512x_xop_1277 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_251_inst
    process(add74_247, shr_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_247, shr_235, tmp_var);
      add79_252 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_448_inst
    process(shr_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_235, type_cast_447_wire_constant, tmp_var);
      tmp554x_xop_449 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_655_inst
    process(tmp540_644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp540_644, type_cast_654_wire_constant, tmp_var);
      tmp540x_xop_656 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_899_inst
    process(tmp524_888) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp524_888, type_cast_898_wire_constant, tmp_var);
      tmp524x_xop_900 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1286_inst
    process(iNsTr_186_1281) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_186_1281, type_cast_1285_wire_constant, tmp_var);
      xx_xop_1287 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1418_inst
    process(indvar_1297) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1297, type_cast_1417_wire_constant, tmp_var);
      indvarx_xnext_1419 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_458_inst
    process(iNsTr_26_453) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_453, type_cast_457_wire_constant, tmp_var);
      xx_xop563_459 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_625_inst
    process(indvar547_469) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar547_469, type_cast_624_wire_constant, tmp_var);
      indvarx_xnext548_626 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_665_inst
    process(iNsTr_39_660) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_660, type_cast_664_wire_constant, tmp_var);
      xx_xop562_666 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_832_inst
    process(indvar531_676) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar531_676, type_cast_831_wire_constant, tmp_var);
      indvarx_xnext532_833 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_909_inst
    process(iNsTr_53_904) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_904, type_cast_908_wire_constant, tmp_var);
      xx_xop561_910 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_944_inst
    process(indvar517_920) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar517_920, type_cast_943_wire_constant, tmp_var);
      indvarx_xnext518_945 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_246_inst
    process(iNsTr_14_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_241, type_cast_245_wire_constant, tmp_var);
      add74_247 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1423_inst
    process(indvarx_xnext_1419, tmp516_1294) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1419, tmp516_1294, tmp_var);
      exitcond1_1424 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_630_inst
    process(indvarx_xnext548_626, tmp559_466) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext548_626, tmp559_466, tmp_var);
      exitcond3_631 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_837_inst
    process(indvarx_xnext532_833, tmp545_673) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext532_833, tmp545_673, tmp_var);
      exitcond2_838 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_949_inst
    process(indvarx_xnext518_945, tmp529_917) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext518_945, tmp529_917, tmp_var);
      exitcond_950 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1044_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_1043_wire_constant, tmp_var);
      shr304_1045 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1100_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_1099_wire_constant, tmp_var);
      shr321_1101 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1156_inst
    process(add79_252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_252, type_cast_1155_wire_constant, tmp_var);
      shr338_1157 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1264_inst
    process(mul259_869) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_869, type_cast_1263_wire_constant, tmp_var);
      tmp512_1265 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_234_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_233_wire_constant, tmp_var);
      shr_235 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_240_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_229, type_cast_239_wire_constant, tmp_var);
      iNsTr_14_241 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_643_inst
    process(mul91_283) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_283, type_cast_642_wire_constant, tmp_var);
      tmp540_644 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_887_inst
    process(mul259_869) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_869, type_cast_886_wire_constant, tmp_var);
      tmp524_888 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1214_inst
    process(sub_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1205, type_cast_1213_wire_constant, tmp_var);
      shr364_1215 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1224_inst
    process(sub_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1205, type_cast_1223_wire_constant, tmp_var);
      shr370_1225 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1234_inst
    process(sub_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1205, type_cast_1233_wire_constant, tmp_var);
      shr376_1235 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1324_inst
    process(tmp425_1315) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp425_1315, type_cast_1323_wire_constant, tmp_var);
      shr432_1325 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1334_inst
    process(tmp425_1315) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp425_1315, type_cast_1333_wire_constant, tmp_var);
      shr438_1335 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1344_inst
    process(tmp425_1315) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp425_1315, type_cast_1343_wire_constant, tmp_var);
      shr444_1345 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1354_inst
    process(tmp425_1315) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp425_1315, type_cast_1353_wire_constant, tmp_var);
      shr450_1355 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1364_inst
    process(tmp425_1315) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp425_1315, type_cast_1363_wire_constant, tmp_var);
      shr456_1365 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1374_inst
    process(tmp425_1315) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp425_1315, type_cast_1373_wire_constant, tmp_var);
      shr462_1375 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1384_inst
    process(tmp425_1315) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp425_1315, type_cast_1383_wire_constant, tmp_var);
      shr468_1385 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_223_inst
    process(conv63_215, conv61_211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_215, conv61_211, tmp_var);
      mul_224 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_228_inst
    process(mul_224, conv65_219) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_224, conv65_219, tmp_var);
      mul66_229 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_272_inst
    process(conv84_260, conv82_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_260, conv82_256, tmp_var);
      mul85_273 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_277_inst
    process(mul85_273, conv87_264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_273, conv87_264, tmp_var);
      mul88_278 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_282_inst
    process(mul88_278, conv90_268) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_278, conv90_268, tmp_var);
      mul91_283 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_863_inst
    process(conv255_855, conv253_851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_855, conv253_851, tmp_var);
      mul256_864 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_868_inst
    process(mul256_864, conv258_859) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_864, conv258_859, tmp_var);
      mul259_869 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_106_inst
    process(shl18_95, conv20_102) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_95, conv20_102, tmp_var);
      add21_107 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_131_inst
    process(shl27_120, conv29_127) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_120, conv29_127, tmp_var);
      add30_132 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_156_inst
    process(shl36_145, conv38_152) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_145, conv38_152, tmp_var);
      add39_157 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_181_inst
    process(shl45_170, conv47_177) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_170, conv47_177, tmp_var);
      add48_182 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_206_inst
    process(shl54_195, conv56_202) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_195, conv56_202, tmp_var);
      add57_207 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_307_inst
    process(shl96_296, conv98_303) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_296, conv98_303, tmp_var);
      add99_308 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_332_inst
    process(shl105_321, conv107_328) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_321, conv107_328, tmp_var);
      add108_333 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_357_inst
    process(shl114_346, conv116_353) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_346, conv116_353, tmp_var);
      add117_358 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_382_inst
    process(shl123_371, conv125_378) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_371, conv125_378, tmp_var);
      add126_383 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_407_inst
    process(shl132_396, conv134_403) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_396, conv134_403, tmp_var);
      add135_408 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_56_inst
    process(shl_45, conv3_52) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_45, conv3_52, tmp_var);
      add_57 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_81_inst
    process(shl9_70, conv11_77) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_70, conv11_77, tmp_var);
      add12_82 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_507_inst
    process(shl146_496, conv149_503) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_496, conv149_503, tmp_var);
      add150_508 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_525_inst
    process(shl152_514, conv155_521) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_514, conv155_521, tmp_var);
      add156_526 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_543_inst
    process(shl158_532, conv161_539) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_532, conv161_539, tmp_var);
      add162_544 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_561_inst
    process(shl164_550, conv167_557) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_550, conv167_557, tmp_var);
      add168_562 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_579_inst
    process(shl170_568, conv173_575) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_568, conv173_575, tmp_var);
      add174_580 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_597_inst
    process(shl176_586, conv179_593) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_586, conv179_593, tmp_var);
      add180_598 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_615_inst
    process(shl182_604, conv185_611) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_604, conv185_611, tmp_var);
      add186_616 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_714_inst
    process(shl202_703, conv205_710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_703, conv205_710, tmp_var);
      add206_715 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_732_inst
    process(shl208_721, conv211_728) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_721, conv211_728, tmp_var);
      add212_733 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_750_inst
    process(shl214_739, conv217_746) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_739, conv217_746, tmp_var);
      add218_751 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_768_inst
    process(shl220_757, conv223_764) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_757, conv223_764, tmp_var);
      add224_769 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_786_inst
    process(shl226_775, conv229_782) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_775, conv229_782, tmp_var);
      add230_787 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_804_inst
    process(shl232_793, conv235_800) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_793, conv235_800, tmp_var);
      add236_805 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_822_inst
    process(shl238_811, conv241_818) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_811, conv241_818, tmp_var);
      add242_823 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_119_inst
    process(conv26_114) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_114, type_cast_118_wire_constant, tmp_var);
      shl27_120 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_144_inst
    process(conv35_139) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_139, type_cast_143_wire_constant, tmp_var);
      shl36_145 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_169_inst
    process(conv44_164) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_164, type_cast_168_wire_constant, tmp_var);
      shl45_170 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_194_inst
    process(conv53_189) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_189, type_cast_193_wire_constant, tmp_var);
      shl54_195 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_295_inst
    process(conv95_290) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_290, type_cast_294_wire_constant, tmp_var);
      shl96_296 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_320_inst
    process(conv104_315) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_315, type_cast_319_wire_constant, tmp_var);
      shl105_321 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_345_inst
    process(conv113_340) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_340, type_cast_344_wire_constant, tmp_var);
      shl114_346 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_370_inst
    process(conv122_365) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_365, type_cast_369_wire_constant, tmp_var);
      shl123_371 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_395_inst
    process(conv131_390) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_390, type_cast_394_wire_constant, tmp_var);
      shl132_396 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_44_inst
    process(conv1_39) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_39, type_cast_43_wire_constant, tmp_var);
      shl_45 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_69_inst
    process(conv8_64) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_64, type_cast_68_wire_constant, tmp_var);
      shl9_70 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_94_inst
    process(conv17_89) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_89, type_cast_93_wire_constant, tmp_var);
      shl18_95 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_495_inst
    process(conv144_490) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_490, type_cast_494_wire_constant, tmp_var);
      shl146_496 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_513_inst
    process(add150_508) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_508, type_cast_512_wire_constant, tmp_var);
      shl152_514 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_531_inst
    process(add156_526) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_526, type_cast_530_wire_constant, tmp_var);
      shl158_532 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_549_inst
    process(add162_544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_544, type_cast_548_wire_constant, tmp_var);
      shl164_550 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_567_inst
    process(add168_562) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_562, type_cast_566_wire_constant, tmp_var);
      shl170_568 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_585_inst
    process(add174_580) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_580, type_cast_584_wire_constant, tmp_var);
      shl176_586 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_603_inst
    process(add180_598) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_598, type_cast_602_wire_constant, tmp_var);
      shl182_604 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_702_inst
    process(conv200_697) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_697, type_cast_701_wire_constant, tmp_var);
      shl202_703 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_720_inst
    process(add206_715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_715, type_cast_719_wire_constant, tmp_var);
      shl208_721 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_738_inst
    process(add212_733) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_733, type_cast_737_wire_constant, tmp_var);
      shl214_739 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_756_inst
    process(add218_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_751, type_cast_755_wire_constant, tmp_var);
      shl220_757 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_774_inst
    process(add224_769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_769, type_cast_773_wire_constant, tmp_var);
      shl226_775 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_792_inst
    process(add230_787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_787, type_cast_791_wire_constant, tmp_var);
      shl232_793 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_810_inst
    process(add236_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_805, type_cast_809_wire_constant, tmp_var);
      shl238_811 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1204_inst
    process(conv355_1200, conv276_968) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv355_1200, conv276_968, tmp_var);
      sub_1205 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1270_inst
    process(tmp512_1265) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp512_1265, type_cast_1269_wire_constant, tmp_var);
      tmp513_1271 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_413_inst
    process(mul66_229) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_229, type_cast_412_wire_constant, tmp_var);
      cmp505_415 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_429_inst
    process(mul91_283) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_283, type_cast_428_wire_constant, tmp_var);
      cmp194501_430 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_442_inst
    process(shr_235) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_235, type_cast_441_wire_constant, tmp_var);
      tmp555_443 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_649_inst
    process(tmp540_644) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp540_644, type_cast_648_wire_constant, tmp_var);
      tmp541_650 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_874_inst
    process(mul259_869) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_869, type_cast_873_wire_constant, tmp_var);
      cmp264497_875 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_893_inst
    process(tmp524_888) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp524_888, type_cast_892_wire_constant, tmp_var);
      tmp525_894 <= tmp_var; --
    end process;
    -- shared split operator group (103) : array_obj_ref_1309_index_offset 
    ApIntAdd_group_103: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1308_scaled;
      array_obj_ref_1309_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1309_index_offset_req_0;
      array_obj_ref_1309_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1309_index_offset_req_1;
      array_obj_ref_1309_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_103_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_103_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_103",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 103
    -- shared split operator group (104) : array_obj_ref_481_index_offset 
    ApIntAdd_group_104: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar547_480_scaled;
      array_obj_ref_481_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_481_index_offset_req_0;
      array_obj_ref_481_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_481_index_offset_req_1;
      array_obj_ref_481_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_104_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_104_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_104",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 104
    -- shared split operator group (105) : array_obj_ref_688_index_offset 
    ApIntAdd_group_105: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar531_687_scaled;
      array_obj_ref_688_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_688_index_offset_req_0;
      array_obj_ref_688_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_688_index_offset_req_1;
      array_obj_ref_688_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_105_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_105_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_105",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 105
    -- shared split operator group (106) : array_obj_ref_932_index_offset 
    ApIntAdd_group_106: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar517_931_scaled;
      array_obj_ref_932_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_932_index_offset_req_0;
      array_obj_ref_932_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_932_index_offset_req_1;
      array_obj_ref_932_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_106_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_106_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_106",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 106
    -- unary operator type_cast_1198_inst
    process(call354_1195) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call354_1195, tmp_var);
      type_cast_1198_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_966_inst
    process(call275_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_962, tmp_var);
      type_cast_966_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1314_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1314_load_0_req_0;
      ptr_deref_1314_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1314_load_0_req_1;
      ptr_deref_1314_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1314_word_address_0;
      ptr_deref_1314_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_618_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_618_store_0_req_0;
      ptr_deref_618_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_618_store_0_req_1;
      ptr_deref_618_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_618_word_address_0;
      data_in <= ptr_deref_618_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_825_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_825_store_0_req_0;
      ptr_deref_825_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_825_store_0_req_1;
      ptr_deref_825_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_825_word_address_0;
      data_in <= ptr_deref_825_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_936_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_936_store_0_req_0;
      ptr_deref_936_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_936_store_0_req_1;
      ptr_deref_936_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_936_word_address_0;
      data_in <= ptr_deref_936_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1182_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1182_inst_req_0;
      RPIPE_Block0_done_1182_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1182_inst_req_1;
      RPIPE_Block0_done_1182_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call346_1183 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1185_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1185_inst_req_0;
      RPIPE_Block1_done_1185_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1185_inst_req_1;
      RPIPE_Block1_done_1185_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call348_1186 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1188_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1188_inst_req_0;
      RPIPE_Block2_done_1188_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1188_inst_req_1;
      RPIPE_Block2_done_1188_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call350_1189 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1191_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1191_inst_req_0;
      RPIPE_Block3_done_1191_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1191_inst_req_1;
      RPIPE_Block3_done_1191_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call352_1192 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_147_inst RPIPE_ConvTranspose_input_pipe_159_inst RPIPE_ConvTranspose_input_pipe_310_inst RPIPE_ConvTranspose_input_pipe_172_inst RPIPE_ConvTranspose_input_pipe_184_inst RPIPE_ConvTranspose_input_pipe_197_inst RPIPE_ConvTranspose_input_pipe_298_inst RPIPE_ConvTranspose_input_pipe_285_inst RPIPE_ConvTranspose_input_pipe_34_inst RPIPE_ConvTranspose_input_pipe_47_inst RPIPE_ConvTranspose_input_pipe_59_inst RPIPE_ConvTranspose_input_pipe_72_inst RPIPE_ConvTranspose_input_pipe_84_inst RPIPE_ConvTranspose_input_pipe_97_inst RPIPE_ConvTranspose_input_pipe_109_inst RPIPE_ConvTranspose_input_pipe_122_inst RPIPE_ConvTranspose_input_pipe_134_inst RPIPE_ConvTranspose_input_pipe_323_inst RPIPE_ConvTranspose_input_pipe_335_inst RPIPE_ConvTranspose_input_pipe_348_inst RPIPE_ConvTranspose_input_pipe_360_inst RPIPE_ConvTranspose_input_pipe_373_inst RPIPE_ConvTranspose_input_pipe_385_inst RPIPE_ConvTranspose_input_pipe_398_inst RPIPE_ConvTranspose_input_pipe_485_inst RPIPE_ConvTranspose_input_pipe_498_inst RPIPE_ConvTranspose_input_pipe_516_inst RPIPE_ConvTranspose_input_pipe_534_inst RPIPE_ConvTranspose_input_pipe_552_inst RPIPE_ConvTranspose_input_pipe_570_inst RPIPE_ConvTranspose_input_pipe_588_inst RPIPE_ConvTranspose_input_pipe_606_inst RPIPE_ConvTranspose_input_pipe_692_inst RPIPE_ConvTranspose_input_pipe_705_inst RPIPE_ConvTranspose_input_pipe_723_inst RPIPE_ConvTranspose_input_pipe_741_inst RPIPE_ConvTranspose_input_pipe_759_inst RPIPE_ConvTranspose_input_pipe_777_inst RPIPE_ConvTranspose_input_pipe_795_inst RPIPE_ConvTranspose_input_pipe_813_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_310_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_298_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_285_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_323_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_335_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_348_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_360_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_373_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_385_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_398_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_485_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_498_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_516_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_534_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_552_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_570_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_588_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_606_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_692_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_705_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_723_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_741_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_759_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_777_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_795_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_813_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_310_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_298_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_285_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_323_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_335_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_348_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_360_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_373_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_385_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_398_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_485_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_498_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_516_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_534_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_552_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_570_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_588_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_606_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_692_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_705_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_723_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_741_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_759_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_777_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_795_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_813_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_310_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_298_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_285_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_323_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_335_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_348_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_360_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_373_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_385_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_398_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_485_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_498_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_516_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_534_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_552_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_570_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_588_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_606_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_692_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_705_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_723_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_741_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_759_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_777_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_795_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_813_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_310_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_298_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_285_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_323_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_335_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_348_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_360_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_373_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_385_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_398_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_485_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_498_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_516_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_534_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_552_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_570_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_588_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_606_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_692_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_705_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_723_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_741_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_759_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_777_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_795_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_813_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call37_148 <= data_out(319 downto 312);
      call41_160 <= data_out(311 downto 304);
      call101_311 <= data_out(303 downto 296);
      call46_173 <= data_out(295 downto 288);
      call50_185 <= data_out(287 downto 280);
      call55_198 <= data_out(279 downto 272);
      call97_299 <= data_out(271 downto 264);
      call92_286 <= data_out(263 downto 256);
      call_35 <= data_out(255 downto 248);
      call2_48 <= data_out(247 downto 240);
      call5_60 <= data_out(239 downto 232);
      call10_73 <= data_out(231 downto 224);
      call14_85 <= data_out(223 downto 216);
      call19_98 <= data_out(215 downto 208);
      call23_110 <= data_out(207 downto 200);
      call28_123 <= data_out(199 downto 192);
      call32_135 <= data_out(191 downto 184);
      call106_324 <= data_out(183 downto 176);
      call110_336 <= data_out(175 downto 168);
      call115_349 <= data_out(167 downto 160);
      call119_361 <= data_out(159 downto 152);
      call124_374 <= data_out(151 downto 144);
      call128_386 <= data_out(143 downto 136);
      call133_399 <= data_out(135 downto 128);
      call143_486 <= data_out(127 downto 120);
      call147_499 <= data_out(119 downto 112);
      call153_517 <= data_out(111 downto 104);
      call159_535 <= data_out(103 downto 96);
      call165_553 <= data_out(95 downto 88);
      call171_571 <= data_out(87 downto 80);
      call177_589 <= data_out(79 downto 72);
      call183_607 <= data_out(71 downto 64);
      call199_693 <= data_out(63 downto 56);
      call203_706 <= data_out(55 downto 48);
      call209_724 <= data_out(47 downto 40);
      call215_742 <= data_out(39 downto 32);
      call221_760 <= data_out(31 downto 24);
      call227_778 <= data_out(23 downto 16);
      call233_796 <= data_out(15 downto 8);
      call239_814 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_1000_inst WPIPE_Block0_start_1004_inst WPIPE_Block0_start_1007_inst WPIPE_Block0_start_1010_inst WPIPE_Block0_start_969_inst WPIPE_Block0_start_972_inst WPIPE_Block0_start_975_inst WPIPE_Block0_start_978_inst WPIPE_Block0_start_981_inst WPIPE_Block0_start_984_inst WPIPE_Block0_start_987_inst WPIPE_Block0_start_990_inst WPIPE_Block0_start_993_inst WPIPE_Block0_start_996_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_1000_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_1004_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_1007_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_1010_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_969_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_972_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_975_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_978_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_981_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_984_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_987_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_990_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_993_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_996_inst_req_0;
      WPIPE_Block0_start_1000_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_1004_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_1007_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_1010_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_969_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_972_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_975_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_978_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_981_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_984_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_987_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_990_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_993_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_996_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_1000_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_1004_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_1007_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_1010_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_969_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_972_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_975_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_978_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_981_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_984_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_987_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_990_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_993_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_996_inst_req_1;
      WPIPE_Block0_start_1000_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_1004_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_1007_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_1010_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_969_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_972_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_975_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_978_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_981_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_984_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_987_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_990_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_993_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_996_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= type_cast_1002_wire_constant & add117_358 & add126_383 & add135_408 & add_57 & add12_82 & add21_107 & add30_132 & add39_157 & add48_182 & add57_207 & add99_308 & add108_333 & type_cast_998_wire_constant;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1031_inst WPIPE_Block1_start_1034_inst WPIPE_Block1_start_1037_inst WPIPE_Block1_start_1050_inst WPIPE_Block1_start_1057_inst WPIPE_Block1_start_1060_inst WPIPE_Block1_start_1063_inst WPIPE_Block1_start_1066_inst WPIPE_Block1_start_1013_inst WPIPE_Block1_start_1016_inst WPIPE_Block1_start_1019_inst WPIPE_Block1_start_1022_inst WPIPE_Block1_start_1025_inst WPIPE_Block1_start_1028_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block1_start_1031_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1034_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1037_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1050_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1057_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1060_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1063_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1066_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1013_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1016_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1019_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1022_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1025_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1028_inst_req_0;
      WPIPE_Block1_start_1031_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1034_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1037_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1050_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1057_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1060_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1063_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1066_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1013_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1016_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1019_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1022_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1025_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1028_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block1_start_1031_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1034_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1037_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1050_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1057_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1060_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1063_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1066_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1013_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1016_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1019_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1022_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1025_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1028_inst_req_1;
      WPIPE_Block1_start_1031_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1034_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1037_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1050_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1057_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1060_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1063_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1066_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1013_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1016_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1019_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1022_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1025_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1028_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add57_207 & add99_308 & add108_333 & conv305_1049 & conv307_1056 & add117_358 & add126_383 & add135_408 & add_57 & add12_82 & add21_107 & add30_132 & add39_157 & add48_182;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1113_inst WPIPE_Block2_start_1116_inst WPIPE_Block2_start_1119_inst WPIPE_Block2_start_1069_inst WPIPE_Block2_start_1072_inst WPIPE_Block2_start_1122_inst WPIPE_Block2_start_1075_inst WPIPE_Block2_start_1078_inst WPIPE_Block2_start_1081_inst WPIPE_Block2_start_1084_inst WPIPE_Block2_start_1087_inst WPIPE_Block2_start_1090_inst WPIPE_Block2_start_1093_inst WPIPE_Block2_start_1106_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block2_start_1113_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1116_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1119_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1069_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1072_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1122_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1075_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1078_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1081_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1084_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1087_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1090_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1093_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1106_inst_req_0;
      WPIPE_Block2_start_1113_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1116_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1119_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1069_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1072_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1122_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1075_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1078_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1081_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1084_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1087_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1090_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1093_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1106_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block2_start_1113_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1116_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1119_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1069_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1072_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1122_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1075_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1078_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1081_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1084_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1087_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1090_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1093_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1106_inst_req_1;
      WPIPE_Block2_start_1113_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1116_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1119_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1069_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1072_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1122_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1075_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1078_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1081_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1084_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1087_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1090_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1093_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1106_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= conv324_1112 & add117_358 & add126_383 & add_57 & add12_82 & add135_408 & add21_107 & add30_132 & add39_157 & add48_182 & add57_207 & add99_308 & add108_333 & conv322_1105;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1149_inst WPIPE_Block3_start_1162_inst WPIPE_Block3_start_1169_inst WPIPE_Block3_start_1172_inst WPIPE_Block3_start_1175_inst WPIPE_Block3_start_1178_inst WPIPE_Block3_start_1125_inst WPIPE_Block3_start_1128_inst WPIPE_Block3_start_1131_inst WPIPE_Block3_start_1134_inst WPIPE_Block3_start_1137_inst WPIPE_Block3_start_1140_inst WPIPE_Block3_start_1143_inst WPIPE_Block3_start_1146_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block3_start_1149_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1162_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1169_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1172_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1175_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1178_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1125_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1128_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1131_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1134_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1137_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1140_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1143_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1146_inst_req_0;
      WPIPE_Block3_start_1149_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1162_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1169_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1172_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1175_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1178_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1125_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1128_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1131_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1134_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1137_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1140_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1143_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1146_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block3_start_1149_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1162_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1169_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1172_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1175_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1178_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1125_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1128_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1131_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1134_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1137_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1140_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1143_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1146_inst_req_1;
      WPIPE_Block3_start_1149_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1162_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1169_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1172_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1175_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1178_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1125_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1128_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1131_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1134_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1137_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1140_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1143_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1146_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add108_333 & conv339_1161 & conv341_1168 & add117_358 & add126_383 & add135_408 & add_57 & add12_82 & add21_107 & add30_132 & add39_157 & add48_182 & add57_207 & add99_308;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1396_inst WPIPE_ConvTranspose_output_pipe_1399_inst WPIPE_ConvTranspose_output_pipe_1402_inst WPIPE_ConvTranspose_output_pipe_1240_inst WPIPE_ConvTranspose_output_pipe_1243_inst WPIPE_ConvTranspose_output_pipe_1405_inst WPIPE_ConvTranspose_output_pipe_1246_inst WPIPE_ConvTranspose_output_pipe_1390_inst WPIPE_ConvTranspose_output_pipe_1249_inst WPIPE_ConvTranspose_output_pipe_1408_inst WPIPE_ConvTranspose_output_pipe_1393_inst WPIPE_ConvTranspose_output_pipe_1411_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal sample_req, sample_ack : BooleanArray( 11 downto 0);
      signal update_req, update_ack : BooleanArray( 11 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 11 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant inBUFs : IntegerArray(11 downto 0) := (11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1396_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1399_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1402_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1240_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1243_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1405_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1246_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1390_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1249_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1408_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1393_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1411_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1396_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1399_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1402_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1240_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1243_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1405_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1246_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1390_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1249_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1408_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1393_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1411_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1396_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1399_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1402_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1240_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1243_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1405_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1246_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1390_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1249_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1408_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1393_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1411_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1396_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1399_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1402_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1240_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1243_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1405_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1246_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1390_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1249_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1408_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1393_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1411_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      data_in <= conv459_1369 & conv453_1359 & conv447_1349 & conv379_1239 & conv373_1229 & conv441_1339 & conv367_1219 & conv471_1389 & conv361_1209 & conv435_1329 & conv465_1379 & conv429_1319;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 12, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_962_call call_stmt_1195_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_962_call_req_0;
      reqL_unguarded(0) <= call_stmt_1195_call_req_0;
      call_stmt_962_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1195_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_962_call_req_1;
      reqR_unguarded(0) <= call_stmt_1195_call_req_1;
      call_stmt_962_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1195_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call275_962 <= data_out(127 downto 64);
      call354_1195 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3646_start: Boolean;
  signal convTransposeA_CP_3646_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1530_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1456_inst_ack_0 : boolean;
  signal type_cast_1538_inst_req_0 : boolean;
  signal type_cast_1538_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1468_inst_ack_0 : boolean;
  signal type_cast_1472_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1459_inst_ack_0 : boolean;
  signal type_cast_1526_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1447_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1468_inst_req_0 : boolean;
  signal type_cast_1538_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1456_inst_req_1 : boolean;
  signal type_cast_1610_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1481_inst_req_0 : boolean;
  signal type_cast_1526_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1456_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1447_inst_req_0 : boolean;
  signal type_cast_1614_inst_ack_1 : boolean;
  signal type_cast_1538_inst_ack_1 : boolean;
  signal type_cast_1472_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1444_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1456_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1459_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1459_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1447_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1450_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1459_inst_req_0 : boolean;
  signal type_cast_1534_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1453_inst_ack_1 : boolean;
  signal type_cast_1534_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1453_inst_req_1 : boolean;
  signal type_cast_1534_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1453_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1453_inst_req_0 : boolean;
  signal addr_of_1655_final_reg_req_1 : boolean;
  signal addr_of_1655_final_reg_ack_1 : boolean;
  signal RPIPE_Block0_start_1481_inst_ack_0 : boolean;
  signal type_cast_1472_inst_req_1 : boolean;
  signal type_cast_1472_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1444_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1447_inst_ack_1 : boolean;
  signal type_cast_1610_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1444_inst_req_1 : boolean;
  signal type_cast_1526_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1462_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1481_inst_req_1 : boolean;
  signal type_cast_1610_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1481_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1444_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1450_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1462_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1468_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1462_inst_req_1 : boolean;
  signal array_obj_ref_1654_index_offset_req_1 : boolean;
  signal type_cast_1526_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1462_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1468_inst_ack_1 : boolean;
  signal type_cast_1618_inst_ack_0 : boolean;
  signal type_cast_1648_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1441_inst_req_0 : boolean;
  signal type_cast_1614_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1441_inst_ack_0 : boolean;
  signal type_cast_1614_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1450_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1465_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1465_inst_ack_0 : boolean;
  signal type_cast_1485_inst_req_0 : boolean;
  signal type_cast_1618_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1465_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1465_inst_ack_1 : boolean;
  signal type_cast_1648_inst_ack_0 : boolean;
  signal type_cast_1530_inst_req_0 : boolean;
  signal array_obj_ref_1654_index_offset_req_0 : boolean;
  signal type_cast_1648_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1441_inst_req_1 : boolean;
  signal type_cast_1530_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1441_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1450_inst_ack_0 : boolean;
  signal type_cast_1618_inst_ack_1 : boolean;
  signal type_cast_1614_inst_req_1 : boolean;
  signal type_cast_1618_inst_req_0 : boolean;
  signal type_cast_1648_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1499_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1499_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1499_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1499_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1496_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1496_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1496_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1496_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1493_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1493_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1493_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1493_inst_req_0 : boolean;
  signal type_cast_1485_inst_ack_1 : boolean;
  signal type_cast_1485_inst_req_1 : boolean;
  signal type_cast_1485_inst_ack_0 : boolean;
  signal type_cast_1530_inst_ack_1 : boolean;
  signal type_cast_1534_inst_req_0 : boolean;
  signal addr_of_1655_final_reg_req_0 : boolean;
  signal addr_of_1655_final_reg_ack_0 : boolean;
  signal type_cast_1610_inst_req_0 : boolean;
  signal array_obj_ref_1654_index_offset_ack_1 : boolean;
  signal array_obj_ref_1654_index_offset_ack_0 : boolean;
  signal ptr_deref_1659_load_0_req_0 : boolean;
  signal ptr_deref_1659_load_0_ack_0 : boolean;
  signal ptr_deref_1659_load_0_req_1 : boolean;
  signal ptr_deref_1659_load_0_ack_1 : boolean;
  signal array_obj_ref_1677_index_offset_req_0 : boolean;
  signal array_obj_ref_1677_index_offset_ack_0 : boolean;
  signal array_obj_ref_1677_index_offset_req_1 : boolean;
  signal array_obj_ref_1677_index_offset_ack_1 : boolean;
  signal addr_of_1678_final_reg_req_0 : boolean;
  signal addr_of_1678_final_reg_ack_0 : boolean;
  signal addr_of_1678_final_reg_req_1 : boolean;
  signal addr_of_1678_final_reg_ack_1 : boolean;
  signal ptr_deref_1681_store_0_req_0 : boolean;
  signal ptr_deref_1681_store_0_ack_0 : boolean;
  signal ptr_deref_1681_store_0_req_1 : boolean;
  signal ptr_deref_1681_store_0_ack_1 : boolean;
  signal type_cast_1686_inst_req_0 : boolean;
  signal type_cast_1686_inst_ack_0 : boolean;
  signal type_cast_1686_inst_req_1 : boolean;
  signal type_cast_1686_inst_ack_1 : boolean;
  signal if_stmt_1699_branch_req_0 : boolean;
  signal if_stmt_1699_branch_ack_1 : boolean;
  signal if_stmt_1699_branch_ack_0 : boolean;
  signal type_cast_1727_inst_req_0 : boolean;
  signal type_cast_1727_inst_ack_0 : boolean;
  signal type_cast_1727_inst_req_1 : boolean;
  signal type_cast_1727_inst_ack_1 : boolean;
  signal type_cast_1743_inst_req_0 : boolean;
  signal type_cast_1743_inst_ack_0 : boolean;
  signal type_cast_1743_inst_req_1 : boolean;
  signal type_cast_1743_inst_ack_1 : boolean;
  signal if_stmt_1750_branch_req_0 : boolean;
  signal if_stmt_1750_branch_ack_1 : boolean;
  signal if_stmt_1750_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1786_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1786_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1786_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1786_inst_ack_1 : boolean;
  signal phi_stmt_1548_req_0 : boolean;
  signal phi_stmt_1555_req_0 : boolean;
  signal phi_stmt_1562_req_0 : boolean;
  signal phi_stmt_1569_req_0 : boolean;
  signal type_cast_1554_inst_req_0 : boolean;
  signal type_cast_1554_inst_ack_0 : boolean;
  signal type_cast_1554_inst_req_1 : boolean;
  signal type_cast_1554_inst_ack_1 : boolean;
  signal phi_stmt_1548_req_1 : boolean;
  signal type_cast_1561_inst_req_0 : boolean;
  signal type_cast_1561_inst_ack_0 : boolean;
  signal type_cast_1561_inst_req_1 : boolean;
  signal type_cast_1561_inst_ack_1 : boolean;
  signal phi_stmt_1555_req_1 : boolean;
  signal type_cast_1568_inst_req_0 : boolean;
  signal type_cast_1568_inst_ack_0 : boolean;
  signal type_cast_1568_inst_req_1 : boolean;
  signal type_cast_1568_inst_ack_1 : boolean;
  signal phi_stmt_1562_req_1 : boolean;
  signal type_cast_1575_inst_req_0 : boolean;
  signal type_cast_1575_inst_ack_0 : boolean;
  signal type_cast_1575_inst_req_1 : boolean;
  signal type_cast_1575_inst_ack_1 : boolean;
  signal phi_stmt_1569_req_1 : boolean;
  signal phi_stmt_1548_ack_0 : boolean;
  signal phi_stmt_1555_ack_0 : boolean;
  signal phi_stmt_1562_ack_0 : boolean;
  signal phi_stmt_1569_ack_0 : boolean;
  signal type_cast_1773_inst_req_0 : boolean;
  signal type_cast_1773_inst_ack_0 : boolean;
  signal type_cast_1773_inst_req_1 : boolean;
  signal type_cast_1773_inst_ack_1 : boolean;
  signal phi_stmt_1770_req_0 : boolean;
  signal phi_stmt_1757_req_1 : boolean;
  signal type_cast_1767_inst_req_0 : boolean;
  signal type_cast_1767_inst_ack_0 : boolean;
  signal type_cast_1767_inst_req_1 : boolean;
  signal type_cast_1767_inst_ack_1 : boolean;
  signal phi_stmt_1764_req_0 : boolean;
  signal type_cast_1775_inst_req_0 : boolean;
  signal type_cast_1775_inst_ack_0 : boolean;
  signal type_cast_1775_inst_req_1 : boolean;
  signal type_cast_1775_inst_ack_1 : boolean;
  signal phi_stmt_1770_req_1 : boolean;
  signal type_cast_1760_inst_req_0 : boolean;
  signal type_cast_1760_inst_ack_0 : boolean;
  signal type_cast_1760_inst_req_1 : boolean;
  signal type_cast_1760_inst_ack_1 : boolean;
  signal phi_stmt_1757_req_0 : boolean;
  signal type_cast_1769_inst_req_0 : boolean;
  signal type_cast_1769_inst_ack_0 : boolean;
  signal type_cast_1769_inst_req_1 : boolean;
  signal type_cast_1769_inst_ack_1 : boolean;
  signal phi_stmt_1764_req_1 : boolean;
  signal phi_stmt_1757_ack_0 : boolean;
  signal phi_stmt_1764_ack_0 : boolean;
  signal phi_stmt_1770_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3646_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3646_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3646_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3646_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3646: Block -- control-path 
    signal convTransposeA_CP_3646_elements: BooleanArray(125 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3646_elements(0) <= convTransposeA_CP_3646_start;
    convTransposeA_CP_3646_symbol <= convTransposeA_CP_3646_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/$entry
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500__entry__
      -- CP-element group 0: 	 branch_block_stmt_1439/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1439/branch_block_stmt_1439__entry__
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_Update/$entry
      -- 
    cr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(0), ack => type_cast_1472_inst_req_1); -- 
    rr_3694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(0), ack => RPIPE_Block0_start_1441_inst_req_0); -- 
    cr_3867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(0), ack => type_cast_1485_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	125 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	84 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1439/assign_stmt_1782__entry__
      -- CP-element group 1: 	 branch_block_stmt_1439/assign_stmt_1782__exit__
      -- CP-element group 1: 	 branch_block_stmt_1439/merge_stmt_1756__exit__
      -- CP-element group 1: 	 branch_block_stmt_1439/assign_stmt_1782/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/assign_stmt_1782/$exit
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/SplitProtocol/Update/cr
      -- 
    rr_4380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(1), ack => type_cast_1554_inst_req_0); -- 
    cr_4385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(1), ack => type_cast_1554_inst_req_1); -- 
    rr_4403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(1), ack => type_cast_1561_inst_req_0); -- 
    cr_4408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(1), ack => type_cast_1561_inst_req_1); -- 
    rr_4426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(1), ack => type_cast_1568_inst_req_0); -- 
    cr_4431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(1), ack => type_cast_1568_inst_req_1); -- 
    rr_4449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(1), ack => type_cast_1575_inst_req_0); -- 
    cr_4454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(1), ack => type_cast_1575_inst_req_1); -- 
    convTransposeA_CP_3646_elements(1) <= convTransposeA_CP_3646_elements(125);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_Update/cr
      -- 
    ra_3695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1441_inst_ack_0, ack => convTransposeA_CP_3646_elements(2)); -- 
    cr_3699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(2), ack => RPIPE_Block0_start_1441_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1441_Update/ca
      -- 
    ca_3700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1441_inst_ack_1, ack => convTransposeA_CP_3646_elements(3)); -- 
    rr_3708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(3), ack => RPIPE_Block0_start_1444_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_Update/cr
      -- 
    ra_3709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1444_inst_ack_0, ack => convTransposeA_CP_3646_elements(4)); -- 
    cr_3713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(4), ack => RPIPE_Block0_start_1444_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1444_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_sample_start_
      -- 
    ca_3714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1444_inst_ack_1, ack => convTransposeA_CP_3646_elements(5)); -- 
    rr_3722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(5), ack => RPIPE_Block0_start_1447_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_update_start_
      -- 
    ra_3723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1447_inst_ack_0, ack => convTransposeA_CP_3646_elements(6)); -- 
    cr_3727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(6), ack => RPIPE_Block0_start_1447_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1447_update_completed_
      -- 
    ca_3728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1447_inst_ack_1, ack => convTransposeA_CP_3646_elements(7)); -- 
    rr_3736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(7), ack => RPIPE_Block0_start_1450_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_Sample/ra
      -- 
    ra_3737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1450_inst_ack_0, ack => convTransposeA_CP_3646_elements(8)); -- 
    cr_3741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(8), ack => RPIPE_Block0_start_1450_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1450_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_Sample/$entry
      -- 
    ca_3742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1450_inst_ack_1, ack => convTransposeA_CP_3646_elements(9)); -- 
    rr_3750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(9), ack => RPIPE_Block0_start_1453_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_update_start_
      -- 
    ra_3751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1453_inst_ack_0, ack => convTransposeA_CP_3646_elements(10)); -- 
    cr_3755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(10), ack => RPIPE_Block0_start_1453_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1453_update_completed_
      -- 
    ca_3756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1453_inst_ack_1, ack => convTransposeA_CP_3646_elements(11)); -- 
    rr_3764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(11), ack => RPIPE_Block0_start_1456_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_sample_completed_
      -- 
    ra_3765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1456_inst_ack_0, ack => convTransposeA_CP_3646_elements(12)); -- 
    cr_3769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(12), ack => RPIPE_Block0_start_1456_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1456_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_Sample/$entry
      -- 
    ca_3770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1456_inst_ack_1, ack => convTransposeA_CP_3646_elements(13)); -- 
    rr_3778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(13), ack => RPIPE_Block0_start_1459_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_update_start_
      -- 
    ra_3779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1459_inst_ack_0, ack => convTransposeA_CP_3646_elements(14)); -- 
    cr_3783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(14), ack => RPIPE_Block0_start_1459_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1459_update_completed_
      -- 
    ca_3784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1459_inst_ack_1, ack => convTransposeA_CP_3646_elements(15)); -- 
    rr_3792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(15), ack => RPIPE_Block0_start_1462_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_Update/cr
      -- 
    ra_3793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1462_inst_ack_0, ack => convTransposeA_CP_3646_elements(16)); -- 
    cr_3797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(16), ack => RPIPE_Block0_start_1462_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1462_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_Sample/rr
      -- 
    ca_3798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1462_inst_ack_1, ack => convTransposeA_CP_3646_elements(17)); -- 
    rr_3806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(17), ack => RPIPE_Block0_start_1465_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_Update/cr
      -- 
    ra_3807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1465_inst_ack_0, ack => convTransposeA_CP_3646_elements(18)); -- 
    cr_3811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(18), ack => RPIPE_Block0_start_1465_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1465_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_sample_start_
      -- 
    ca_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1465_inst_ack_1, ack => convTransposeA_CP_3646_elements(19)); -- 
    rr_3820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(19), ack => RPIPE_Block0_start_1468_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_sample_completed_
      -- 
    ra_3821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1468_inst_ack_0, ack => convTransposeA_CP_3646_elements(20)); -- 
    cr_3825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(20), ack => RPIPE_Block0_start_1468_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1468_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_sample_start_
      -- 
    ca_3826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1468_inst_ack_1, ack => convTransposeA_CP_3646_elements(21)); -- 
    rr_3834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(21), ack => type_cast_1472_inst_req_0); -- 
    rr_3848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(21), ack => RPIPE_Block0_start_1481_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_sample_completed_
      -- 
    ra_3835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1472_inst_ack_0, ack => convTransposeA_CP_3646_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1472_update_completed_
      -- 
    ca_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1472_inst_ack_1, ack => convTransposeA_CP_3646_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_update_start_
      -- 
    ra_3849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1481_inst_ack_0, ack => convTransposeA_CP_3646_elements(24)); -- 
    cr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(24), ack => RPIPE_Block0_start_1481_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1481_update_completed_
      -- 
    ca_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1481_inst_ack_1, ack => convTransposeA_CP_3646_elements(25)); -- 
    rr_3862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(25), ack => type_cast_1485_inst_req_0); -- 
    rr_3876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(25), ack => RPIPE_Block0_start_1493_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_Sample/ra
      -- 
    ra_3863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1485_inst_ack_0, ack => convTransposeA_CP_3646_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/type_cast_1485_Update/$exit
      -- 
    ca_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1485_inst_ack_1, ack => convTransposeA_CP_3646_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_sample_completed_
      -- 
    ra_3877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1493_inst_ack_0, ack => convTransposeA_CP_3646_elements(28)); -- 
    cr_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(28), ack => RPIPE_Block0_start_1493_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1493_update_completed_
      -- 
    ca_3882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1493_inst_ack_1, ack => convTransposeA_CP_3646_elements(29)); -- 
    rr_3890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(29), ack => RPIPE_Block0_start_1496_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_sample_completed_
      -- 
    ra_3891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1496_inst_ack_0, ack => convTransposeA_CP_3646_elements(30)); -- 
    cr_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(30), ack => RPIPE_Block0_start_1496_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1496_update_completed_
      -- 
    ca_3896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1496_inst_ack_1, ack => convTransposeA_CP_3646_elements(31)); -- 
    rr_3904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(31), ack => RPIPE_Block0_start_1499_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_sample_completed_
      -- 
    ra_3905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1499_inst_ack_0, ack => convTransposeA_CP_3646_elements(32)); -- 
    cr_3909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(32), ack => RPIPE_Block0_start_1499_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/RPIPE_Block0_start_1499_update_completed_
      -- 
    ca_3910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1499_inst_ack_1, ack => convTransposeA_CP_3646_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545__entry__
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500/$exit
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1442_to_assign_stmt_1500__exit__
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/$entry
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_sample_start_
      -- 
    cr_3940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(34), ack => type_cast_1530_inst_req_1); -- 
    rr_3963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(34), ack => type_cast_1538_inst_req_0); -- 
    cr_3968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(34), ack => type_cast_1538_inst_req_1); -- 
    rr_3921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(34), ack => type_cast_1526_inst_req_0); -- 
    cr_3954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(34), ack => type_cast_1534_inst_req_1); -- 
    cr_3926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(34), ack => type_cast_1526_inst_req_1); -- 
    rr_3935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(34), ack => type_cast_1530_inst_req_0); -- 
    rr_3949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(34), ack => type_cast_1534_inst_req_0); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(23) & convTransposeA_CP_3646_elements(27) & convTransposeA_CP_3646_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_sample_completed_
      -- 
    ra_3922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1526_inst_ack_0, ack => convTransposeA_CP_3646_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1526_update_completed_
      -- 
    ca_3927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1526_inst_ack_1, ack => convTransposeA_CP_3646_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_Sample/ra
      -- 
    ra_3936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1530_inst_ack_0, ack => convTransposeA_CP_3646_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1530_Update/ca
      -- 
    ca_3941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1530_inst_ack_1, ack => convTransposeA_CP_3646_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_sample_completed_
      -- 
    ra_3950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1534_inst_ack_0, ack => convTransposeA_CP_3646_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1534_Update/$exit
      -- 
    ca_3955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1534_inst_ack_1, ack => convTransposeA_CP_3646_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_Sample/$exit
      -- 
    ra_3964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1538_inst_ack_0, ack => convTransposeA_CP_3646_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/type_cast_1538_Update/ca
      -- 
    ca_3969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1538_inst_ack_1, ack => convTransposeA_CP_3646_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1439/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545__exit__
      -- CP-element group 43: 	 branch_block_stmt_1439/assign_stmt_1507_to_assign_stmt_1545/$exit
      -- CP-element group 43: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1548/$entry
      -- CP-element group 43: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1555/$entry
      -- CP-element group 43: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1562/$entry
      -- CP-element group 43: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1569/$entry
      -- CP-element group 43: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/$entry
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(36) & convTransposeA_CP_3646_elements(38) & convTransposeA_CP_3646_elements(40) & convTransposeA_CP_3646_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	102 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_sample_completed_
      -- 
    ra_3981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1610_inst_ack_0, ack => convTransposeA_CP_3646_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	102 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_Update/ca
      -- 
    ca_3986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1610_inst_ack_1, ack => convTransposeA_CP_3646_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	102 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_Sample/ra
      -- 
    ra_3995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1614_inst_ack_0, ack => convTransposeA_CP_3646_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	102 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_update_completed_
      -- 
    ca_4000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1614_inst_ack_1, ack => convTransposeA_CP_3646_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	102 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_Sample/$exit
      -- 
    ra_4009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1618_inst_ack_0, ack => convTransposeA_CP_3646_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	102 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_Update/ca
      -- 
    ca_4014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1618_inst_ack_1, ack => convTransposeA_CP_3646_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	102 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_Sample/$exit
      -- 
    ra_4023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1648_inst_ack_0, ack => convTransposeA_CP_3646_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	102 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_final_index_sum_regn_Sample/req
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_index_scaled_1
      -- 
    ca_4028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1648_inst_ack_1, ack => convTransposeA_CP_3646_elements(51)); -- 
    req_4053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(51), ack => array_obj_ref_1654_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_final_index_sum_regn_Sample/ack
      -- 
    ack_4054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1654_index_offset_ack_0, ack => convTransposeA_CP_3646_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	102 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_request/req
      -- CP-element group 53: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_final_index_sum_regn_Update/ack
      -- 
    ack_4059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1654_index_offset_ack_1, ack => convTransposeA_CP_3646_elements(53)); -- 
    req_4068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(53), ack => addr_of_1655_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_request/ack
      -- 
    ack_4069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1655_final_reg_ack_0, ack => convTransposeA_CP_3646_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	102 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Sample/word_access_start/word_0/rr
      -- 
    ack_4074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1655_final_reg_ack_1, ack => convTransposeA_CP_3646_elements(55)); -- 
    rr_4107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(55), ack => ptr_deref_1659_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Sample/word_access_start/word_0/ra
      -- 
    ra_4108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1659_load_0_ack_0, ack => convTransposeA_CP_3646_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	102 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/ptr_deref_1659_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/ptr_deref_1659_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/ptr_deref_1659_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/ptr_deref_1659_Merge/merge_ack
      -- 
    ca_4119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1659_load_0_ack_1, ack => convTransposeA_CP_3646_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_final_index_sum_regn_Sample/req
      -- 
    req_4149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(58), ack => array_obj_ref_1677_index_offset_req_0); -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(45) & convTransposeA_CP_3646_elements(47) & convTransposeA_CP_3646_elements(49);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_final_index_sum_regn_Sample/ack
      -- 
    ack_4150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1677_index_offset_ack_0, ack => convTransposeA_CP_3646_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	102 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_request/req
      -- 
    ack_4155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1677_index_offset_ack_1, ack => convTransposeA_CP_3646_elements(60)); -- 
    req_4164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(60), ack => addr_of_1678_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_request/ack
      -- 
    ack_4165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1678_final_reg_ack_0, ack => convTransposeA_CP_3646_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	102 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_word_addrgen/root_register_ack
      -- 
    ack_4170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1678_final_reg_ack_1, ack => convTransposeA_CP_3646_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/ptr_deref_1681_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/ptr_deref_1681_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/ptr_deref_1681_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/ptr_deref_1681_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/word_access_start/word_0/rr
      -- 
    rr_4208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(63), ack => ptr_deref_1681_store_0_req_0); -- 
    convTransposeA_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(57) & convTransposeA_CP_3646_elements(62);
      gj_convTransposeA_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Sample/word_access_start/word_0/ra
      -- 
    ra_4209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1681_store_0_ack_0, ack => convTransposeA_CP_3646_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	102 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Update/word_access_complete/word_0/ca
      -- 
    ca_4220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1681_store_0_ack_1, ack => convTransposeA_CP_3646_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_Sample/ra
      -- 
    ra_4229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1686_inst_ack_0, ack => convTransposeA_CP_3646_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	102 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_Update/ca
      -- 
    ca_4234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1686_inst_ack_1, ack => convTransposeA_CP_3646_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698__exit__
      -- CP-element group 68: 	 branch_block_stmt_1439/if_stmt_1699__entry__
      -- CP-element group 68: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/$exit
      -- CP-element group 68: 	 branch_block_stmt_1439/if_stmt_1699_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1439/if_stmt_1699_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1439/if_stmt_1699_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1439/if_stmt_1699_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1439/R_cmp_1700_place
      -- CP-element group 68: 	 branch_block_stmt_1439/if_stmt_1699_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1439/if_stmt_1699_else_link/$entry
      -- 
    branch_req_4242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(68), ack => if_stmt_1699_branch_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(52) & convTransposeA_CP_3646_elements(59) & convTransposeA_CP_3646_elements(65) & convTransposeA_CP_3646_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	111 
    -- CP-element group 69: 	112 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	115 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	118 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1439/assign_stmt_1711__entry__
      -- CP-element group 69: 	 branch_block_stmt_1439/merge_stmt_1705__exit__
      -- CP-element group 69: 	 branch_block_stmt_1439/assign_stmt_1711__exit__
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123
      -- CP-element group 69: 	 branch_block_stmt_1439/if_stmt_1699_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1439/if_stmt_1699_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1439/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1439/assign_stmt_1711/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/assign_stmt_1711/$exit
      -- CP-element group 69: 	 branch_block_stmt_1439/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1439/merge_stmt_1705_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1439/merge_stmt_1705_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/merge_stmt_1705_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1439/merge_stmt_1705_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1699_branch_ack_1, ack => convTransposeA_CP_3646_elements(69)); -- 
    rr_4564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(69), ack => type_cast_1775_inst_req_0); -- 
    cr_4569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(69), ack => type_cast_1775_inst_req_1); -- 
    rr_4587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(69), ack => type_cast_1760_inst_req_0); -- 
    cr_4592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(69), ack => type_cast_1760_inst_req_1); -- 
    rr_4610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(69), ack => type_cast_1769_inst_req_0); -- 
    cr_4615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(69), ack => type_cast_1769_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1439/merge_stmt_1713__exit__
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749__entry__
      -- CP-element group 70: 	 branch_block_stmt_1439/if_stmt_1699_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1439/if_stmt_1699_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1439/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/$entry
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1439/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1439/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1439/merge_stmt_1713_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1439/merge_stmt_1713_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1439/merge_stmt_1713_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1439/merge_stmt_1713_PhiAck/dummy
      -- 
    else_choice_transition_4251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1699_branch_ack_0, ack => convTransposeA_CP_3646_elements(70)); -- 
    rr_4267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(70), ack => type_cast_1727_inst_req_0); -- 
    cr_4272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(70), ack => type_cast_1727_inst_req_1); -- 
    cr_4286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(70), ack => type_cast_1743_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_Sample/ra
      -- 
    ra_4268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1727_inst_ack_0, ack => convTransposeA_CP_3646_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1727_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_Sample/rr
      -- 
    ca_4273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1727_inst_ack_1, ack => convTransposeA_CP_3646_elements(72)); -- 
    rr_4281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(72), ack => type_cast_1743_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_Sample/ra
      -- 
    ra_4282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1743_inst_ack_0, ack => convTransposeA_CP_3646_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749__exit__
      -- CP-element group 74: 	 branch_block_stmt_1439/if_stmt_1750__entry__
      -- CP-element group 74: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/$exit
      -- CP-element group 74: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1439/assign_stmt_1719_to_assign_stmt_1749/type_cast_1743_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1439/if_stmt_1750_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1439/if_stmt_1750_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1439/if_stmt_1750_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1439/if_stmt_1750_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1439/R_cmp112_1751_place
      -- CP-element group 74: 	 branch_block_stmt_1439/if_stmt_1750_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1439/if_stmt_1750_else_link/$entry
      -- 
    ca_4287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1743_inst_ack_1, ack => convTransposeA_CP_3646_elements(74)); -- 
    branch_req_4295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(74), ack => if_stmt_1750_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1439/merge_stmt_1784__exit__
      -- CP-element group 75: 	 branch_block_stmt_1439/assign_stmt_1789__entry__
      -- CP-element group 75: 	 branch_block_stmt_1439/if_stmt_1750_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1439/if_stmt_1750_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1439/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1439/assign_stmt_1789/$entry
      -- CP-element group 75: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_1439/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1439/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1439/merge_stmt_1784_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1439/merge_stmt_1784_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1439/merge_stmt_1784_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1439/merge_stmt_1784_PhiAck/dummy
      -- 
    if_choice_transition_4300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1750_branch_ack_1, ack => convTransposeA_CP_3646_elements(75)); -- 
    req_4320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(75), ack => WPIPE_Block0_done_1786_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	103 
    -- CP-element group 76: 	104 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	108 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1439/if_stmt_1750_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1439/if_stmt_1750_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1757/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1750_branch_ack_0, ack => convTransposeA_CP_3646_elements(76)); -- 
    rr_4507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(76), ack => type_cast_1773_inst_req_0); -- 
    cr_4512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(76), ack => type_cast_1773_inst_req_1); -- 
    rr_4538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(76), ack => type_cast_1767_inst_req_0); -- 
    cr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(76), ack => type_cast_1767_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_Update/req
      -- 
    ack_4321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1786_inst_ack_0, ack => convTransposeA_CP_3646_elements(77)); -- 
    req_4325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(77), ack => WPIPE_Block0_done_1786_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1439/$exit
      -- CP-element group 78: 	 branch_block_stmt_1439/assign_stmt_1789__exit__
      -- CP-element group 78: 	 branch_block_stmt_1439/return__
      -- CP-element group 78: 	 branch_block_stmt_1439/merge_stmt_1791__exit__
      -- CP-element group 78: 	 branch_block_stmt_1439/branch_block_stmt_1439__exit__
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1439/assign_stmt_1789/$exit
      -- CP-element group 78: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1439/assign_stmt_1789/WPIPE_Block0_done_1786_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1439/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1439/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1439/merge_stmt_1791_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1439/merge_stmt_1791_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1439/merge_stmt_1791_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1439/merge_stmt_1791_PhiAck/dummy
      -- 
    ack_4326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1786_inst_ack_1, ack => convTransposeA_CP_3646_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1548/$exit
      -- CP-element group 79: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1552_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_req
      -- 
    phi_stmt_1548_req_4337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1548_req_4337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(79), ack => phi_stmt_1548_req_0); -- 
    -- Element group convTransposeA_CP_3646_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3646_elements(43), ack => convTransposeA_CP_3646_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1555/$exit
      -- CP-element group 80: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1559_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_req
      -- 
    phi_stmt_1555_req_4345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1555_req_4345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(80), ack => phi_stmt_1555_req_0); -- 
    -- Element group convTransposeA_CP_3646_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeA_CP_3646_elements(43), ack => convTransposeA_CP_3646_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1562/$exit
      -- CP-element group 81: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1566_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_req
      -- 
    phi_stmt_1562_req_4353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1562_req_4353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(81), ack => phi_stmt_1562_req_0); -- 
    -- Element group convTransposeA_CP_3646_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeA_CP_3646_elements(43), ack => convTransposeA_CP_3646_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1569/$exit
      -- CP-element group 82: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1573_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_req
      -- 
    phi_stmt_1569_req_4361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1569_req_4361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(82), ack => phi_stmt_1569_req_0); -- 
    -- Element group convTransposeA_CP_3646_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeA_CP_3646_elements(43), ack => convTransposeA_CP_3646_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	97 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1439/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(79) & convTransposeA_CP_3646_elements(80) & convTransposeA_CP_3646_elements(81) & convTransposeA_CP_3646_elements(82);
      gj_convTransposeA_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/SplitProtocol/Sample/ra
      -- 
    ra_4381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1554_inst_ack_0, ack => convTransposeA_CP_3646_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/SplitProtocol/Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/SplitProtocol/Update/ca
      -- 
    ca_4386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1554_inst_ack_1, ack => convTransposeA_CP_3646_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	96 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/$exit
      -- CP-element group 86: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/$exit
      -- CP-element group 86: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_sources/type_cast_1554/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1548/phi_stmt_1548_req
      -- 
    phi_stmt_1548_req_4387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1548_req_4387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(86), ack => phi_stmt_1548_req_1); -- 
    convTransposeA_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(84) & convTransposeA_CP_3646_elements(85);
      gj_convTransposeA_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/SplitProtocol/Sample/ra
      -- 
    ra_4404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1561_inst_ack_0, ack => convTransposeA_CP_3646_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/SplitProtocol/Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/SplitProtocol/Update/ca
      -- 
    ca_4409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1561_inst_ack_1, ack => convTransposeA_CP_3646_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/$exit
      -- CP-element group 89: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/$exit
      -- CP-element group 89: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_sources/type_cast_1561/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1555/phi_stmt_1555_req
      -- 
    phi_stmt_1555_req_4410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1555_req_4410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(89), ack => phi_stmt_1555_req_1); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(87) & convTransposeA_CP_3646_elements(88);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/SplitProtocol/Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/SplitProtocol/Sample/ra
      -- 
    ra_4427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1568_inst_ack_0, ack => convTransposeA_CP_3646_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/SplitProtocol/Update/ca
      -- 
    ca_4432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1568_inst_ack_1, ack => convTransposeA_CP_3646_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/$exit
      -- CP-element group 92: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/$exit
      -- CP-element group 92: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_sources/type_cast_1568/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1562/phi_stmt_1562_req
      -- 
    phi_stmt_1562_req_4433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1562_req_4433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(92), ack => phi_stmt_1562_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(90) & convTransposeA_CP_3646_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/SplitProtocol/Sample/ra
      -- 
    ra_4450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1575_inst_ack_0, ack => convTransposeA_CP_3646_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/SplitProtocol/Update/ca
      -- 
    ca_4455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1575_inst_ack_1, ack => convTransposeA_CP_3646_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/$exit
      -- CP-element group 95: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/$exit
      -- CP-element group 95: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_sources/type_cast_1575/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1569/phi_stmt_1569_req
      -- 
    phi_stmt_1569_req_4456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1569_req_4456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(95), ack => phi_stmt_1569_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(93) & convTransposeA_CP_3646_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	86 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1439/ifx_xend123_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(86) & convTransposeA_CP_3646_elements(89) & convTransposeA_CP_3646_elements(92) & convTransposeA_CP_3646_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  merge  fork  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	83 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	100 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1439/merge_stmt_1547_PhiReqMerge
      -- CP-element group 97: 	 branch_block_stmt_1439/merge_stmt_1547_PhiAck/$entry
      -- 
    convTransposeA_CP_3646_elements(97) <= OrReduce(convTransposeA_CP_3646_elements(83) & convTransposeA_CP_3646_elements(96));
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1439/merge_stmt_1547_PhiAck/phi_stmt_1548_ack
      -- 
    phi_stmt_1548_ack_4461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1548_ack_0, ack => convTransposeA_CP_3646_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1439/merge_stmt_1547_PhiAck/phi_stmt_1555_ack
      -- 
    phi_stmt_1555_ack_4462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1555_ack_0, ack => convTransposeA_CP_3646_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1439/merge_stmt_1547_PhiAck/phi_stmt_1562_ack
      -- 
    phi_stmt_1562_ack_4463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1562_ack_0, ack => convTransposeA_CP_3646_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1439/merge_stmt_1547_PhiAck/phi_stmt_1569_ack
      -- 
    phi_stmt_1569_ack_4464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1569_ack_0, ack => convTransposeA_CP_3646_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	44 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	46 
    -- CP-element group 102: 	47 
    -- CP-element group 102: 	48 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	50 
    -- CP-element group 102: 	51 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	55 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	60 
    -- CP-element group 102: 	62 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	66 
    -- CP-element group 102: 	67 
    -- CP-element group 102:  members (56) 
      -- CP-element group 102: 	 branch_block_stmt_1439/merge_stmt_1547__exit__
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698__entry__
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1655_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1614_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1618_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1648_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1610_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1654_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1659_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/array_obj_ref_1677_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/addr_of_1678_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/ptr_deref_1681_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1439/assign_stmt_1582_to_assign_stmt_1698/type_cast_1686_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1439/merge_stmt_1547_PhiAck/$exit
      -- 
    cr_3985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => type_cast_1610_inst_req_1); -- 
    req_4073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => addr_of_1655_final_reg_req_1); -- 
    req_4058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => array_obj_ref_1654_index_offset_req_1); -- 
    rr_4022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => type_cast_1648_inst_req_0); -- 
    rr_3994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => type_cast_1614_inst_req_0); -- 
    cr_4013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => type_cast_1618_inst_req_1); -- 
    cr_3999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => type_cast_1614_inst_req_1); -- 
    rr_4008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => type_cast_1618_inst_req_0); -- 
    cr_4027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => type_cast_1648_inst_req_1); -- 
    rr_3980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => type_cast_1610_inst_req_0); -- 
    cr_4118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => ptr_deref_1659_load_0_req_1); -- 
    req_4154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => array_obj_ref_1677_index_offset_req_1); -- 
    req_4169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => addr_of_1678_final_reg_req_1); -- 
    cr_4219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => ptr_deref_1681_store_0_req_1); -- 
    rr_4228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => type_cast_1686_inst_req_0); -- 
    cr_4233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(102), ack => type_cast_1686_inst_req_1); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(98) & convTransposeA_CP_3646_elements(99) & convTransposeA_CP_3646_elements(100) & convTransposeA_CP_3646_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	76 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Sample/ra
      -- 
    ra_4508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1773_inst_ack_0, ack => convTransposeA_CP_3646_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	76 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Update/ca
      -- 
    ca_4513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1773_inst_ack_1, ack => convTransposeA_CP_3646_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	110 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/$exit
      -- CP-element group 105: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/$exit
      -- CP-element group 105: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/$exit
      -- CP-element group 105: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_req
      -- 
    phi_stmt_1770_req_4514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1770_req_4514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(105), ack => phi_stmt_1770_req_0); -- 
    convTransposeA_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(103) & convTransposeA_CP_3646_elements(104);
      gj_convTransposeA_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  output  delay-element  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	110 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1757/$exit
      -- CP-element group 106: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/$exit
      -- CP-element group 106: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1763_konst_delay_trans
      -- CP-element group 106: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_req
      -- 
    phi_stmt_1757_req_4522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1757_req_4522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(106), ack => phi_stmt_1757_req_1); -- 
    -- Element group convTransposeA_CP_3646_elements(106) is a control-delay.
    cp_element_106_delay: control_delay_element  generic map(name => " 106_delay", delay_value => 1)  port map(req => convTransposeA_CP_3646_elements(76), ack => convTransposeA_CP_3646_elements(106), clk => clk, reset =>reset);
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/SplitProtocol/Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/SplitProtocol/Sample/ra
      -- 
    ra_4539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1767_inst_ack_0, ack => convTransposeA_CP_3646_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/SplitProtocol/Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/SplitProtocol/Update/ca
      -- 
    ca_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1767_inst_ack_1, ack => convTransposeA_CP_3646_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/$exit
      -- CP-element group 109: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/$exit
      -- CP-element group 109: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1767/SplitProtocol/$exit
      -- CP-element group 109: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_req
      -- 
    phi_stmt_1764_req_4545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1764_req_4545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(109), ack => phi_stmt_1764_req_0); -- 
    convTransposeA_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(107) & convTransposeA_CP_3646_elements(108);
      gj_convTransposeA_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	105 
    -- CP-element group 110: 	106 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	121 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1439/ifx_xelse_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(105) & convTransposeA_CP_3646_elements(106) & convTransposeA_CP_3646_elements(109);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	69 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/SplitProtocol/Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/SplitProtocol/Sample/ra
      -- 
    ra_4565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1775_inst_ack_0, ack => convTransposeA_CP_3646_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	69 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/SplitProtocol/Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/SplitProtocol/Update/ca
      -- 
    ca_4570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1775_inst_ack_1, ack => convTransposeA_CP_3646_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/$exit
      -- CP-element group 113: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/$exit
      -- CP-element group 113: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/$exit
      -- CP-element group 113: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1775/SplitProtocol/$exit
      -- CP-element group 113: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1770/phi_stmt_1770_req
      -- 
    phi_stmt_1770_req_4571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1770_req_4571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(113), ack => phi_stmt_1770_req_1); -- 
    convTransposeA_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(111) & convTransposeA_CP_3646_elements(112);
      gj_convTransposeA_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/SplitProtocol/Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/SplitProtocol/Sample/ra
      -- 
    ra_4588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1760_inst_ack_0, ack => convTransposeA_CP_3646_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	69 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/SplitProtocol/Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/SplitProtocol/Update/ca
      -- 
    ca_4593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1760_inst_ack_1, ack => convTransposeA_CP_3646_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	120 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/$exit
      -- CP-element group 116: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/$exit
      -- CP-element group 116: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_sources/type_cast_1760/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1757/phi_stmt_1757_req
      -- 
    phi_stmt_1757_req_4594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1757_req_4594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(116), ack => phi_stmt_1757_req_0); -- 
    convTransposeA_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(114) & convTransposeA_CP_3646_elements(115);
      gj_convTransposeA_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/SplitProtocol/Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/SplitProtocol/Sample/ra
      -- 
    ra_4611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1769_inst_ack_0, ack => convTransposeA_CP_3646_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	69 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/SplitProtocol/Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/SplitProtocol/Update/ca
      -- 
    ca_4616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1769_inst_ack_1, ack => convTransposeA_CP_3646_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/$exit
      -- CP-element group 119: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/$exit
      -- CP-element group 119: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_sources/type_cast_1769/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1764/phi_stmt_1764_req
      -- 
    phi_stmt_1764_req_4617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1764_req_4617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3646_elements(119), ack => phi_stmt_1764_req_1); -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(117) & convTransposeA_CP_3646_elements(118);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1439/ifx_xthen_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(113) & convTransposeA_CP_3646_elements(116) & convTransposeA_CP_3646_elements(119);
      gj_convTransposeA_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	110 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1439/merge_stmt_1756_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_1439/merge_stmt_1756_PhiAck/$entry
      -- 
    convTransposeA_CP_3646_elements(121) <= OrReduce(convTransposeA_CP_3646_elements(110) & convTransposeA_CP_3646_elements(120));
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1439/merge_stmt_1756_PhiAck/phi_stmt_1757_ack
      -- 
    phi_stmt_1757_ack_4622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1757_ack_0, ack => convTransposeA_CP_3646_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1439/merge_stmt_1756_PhiAck/phi_stmt_1764_ack
      -- 
    phi_stmt_1764_ack_4623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1764_ack_0, ack => convTransposeA_CP_3646_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1439/merge_stmt_1756_PhiAck/phi_stmt_1770_ack
      -- 
    phi_stmt_1770_ack_4624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1770_ack_0, ack => convTransposeA_CP_3646_elements(124)); -- 
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	1 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1439/merge_stmt_1756_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3646_elements(122) & convTransposeA_CP_3646_elements(123) & convTransposeA_CP_3646_elements(124);
      gj_convTransposeA_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3646_elements(125), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom81_1676_resized : std_logic_vector(13 downto 0);
    signal R_idxprom81_1676_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1653_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1653_scaled : std_logic_vector(13 downto 0);
    signal add41_1507 : std_logic_vector(15 downto 0);
    signal add54_1518 : std_logic_vector(15 downto 0);
    signal add73_1629 : std_logic_vector(63 downto 0);
    signal add75_1639 : std_logic_vector(63 downto 0);
    signal add86_1693 : std_logic_vector(31 downto 0);
    signal add93_1711 : std_logic_vector(15 downto 0);
    signal add_1491 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1587 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1654_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1654_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1654_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1654_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1654_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1654_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1677_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1677_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1677_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1677_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1677_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1677_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1656 : std_logic_vector(31 downto 0);
    signal arrayidx82_1679 : std_logic_vector(31 downto 0);
    signal call11_1460 : std_logic_vector(15 downto 0);
    signal call13_1463 : std_logic_vector(15 downto 0);
    signal call14_1466 : std_logic_vector(15 downto 0);
    signal call15_1469 : std_logic_vector(15 downto 0);
    signal call16_1482 : std_logic_vector(15 downto 0);
    signal call18_1494 : std_logic_vector(15 downto 0);
    signal call1_1445 : std_logic_vector(15 downto 0);
    signal call20_1497 : std_logic_vector(15 downto 0);
    signal call22_1500 : std_logic_vector(15 downto 0);
    signal call3_1448 : std_logic_vector(15 downto 0);
    signal call5_1451 : std_logic_vector(15 downto 0);
    signal call7_1454 : std_logic_vector(15 downto 0);
    signal call9_1457 : std_logic_vector(15 downto 0);
    signal call_1442 : std_logic_vector(15 downto 0);
    signal cmp101_1724 : std_logic_vector(0 downto 0);
    signal cmp112_1749 : std_logic_vector(0 downto 0);
    signal cmp_1698 : std_logic_vector(0 downto 0);
    signal conv107_1744 : std_logic_vector(31 downto 0);
    signal conv110_1539 : std_logic_vector(31 downto 0);
    signal conv17_1486 : std_logic_vector(31 downto 0);
    signal conv61_1611 : std_logic_vector(63 downto 0);
    signal conv64_1527 : std_logic_vector(63 downto 0);
    signal conv66_1615 : std_logic_vector(63 downto 0);
    signal conv69_1531 : std_logic_vector(63 downto 0);
    signal conv71_1619 : std_logic_vector(63 downto 0);
    signal conv85_1687 : std_logic_vector(31 downto 0);
    signal conv89_1535 : std_logic_vector(31 downto 0);
    signal conv_1473 : std_logic_vector(31 downto 0);
    signal idxprom81_1672 : std_logic_vector(63 downto 0);
    signal idxprom_1649 : std_logic_vector(63 downto 0);
    signal inc105_1728 : std_logic_vector(15 downto 0);
    signal inc105x_xinput_dim0x_x2_1733 : std_logic_vector(15 downto 0);
    signal inc_1719 : std_logic_vector(15 downto 0);
    signal indvar_1548 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1782 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1770 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1569 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1764 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1562 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1740 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1757 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1555 : std_logic_vector(15 downto 0);
    signal mul50_1602 : std_logic_vector(15 downto 0);
    signal mul72_1624 : std_logic_vector(63 downto 0);
    signal mul74_1634 : std_logic_vector(63 downto 0);
    signal mul_1592 : std_logic_vector(15 downto 0);
    signal ptr_deref_1659_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1659_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1659_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1659_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1659_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1681_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1681_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1681_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1681_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1681_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1681_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1479 : std_logic_vector(31 downto 0);
    signal shr111126_1545 : std_logic_vector(31 downto 0);
    signal shr80_1666 : std_logic_vector(63 downto 0);
    signal shr_1645 : std_logic_vector(31 downto 0);
    signal sub44_1597 : std_logic_vector(15 downto 0);
    signal sub57_1523 : std_logic_vector(15 downto 0);
    signal sub58_1607 : std_logic_vector(15 downto 0);
    signal sub_1512 : std_logic_vector(15 downto 0);
    signal tmp1_1582 : std_logic_vector(31 downto 0);
    signal tmp78_1660 : std_logic_vector(63 downto 0);
    signal type_cast_1477_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1505_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1516_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1543_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1552_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1554_wire : std_logic_vector(31 downto 0);
    signal type_cast_1559_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1561_wire : std_logic_vector(15 downto 0);
    signal type_cast_1566_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1568_wire : std_logic_vector(15 downto 0);
    signal type_cast_1573_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1575_wire : std_logic_vector(15 downto 0);
    signal type_cast_1580_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1643_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1664_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1670_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1691_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1709_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1717_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1737_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1760_wire : std_logic_vector(15 downto 0);
    signal type_cast_1763_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1767_wire : std_logic_vector(15 downto 0);
    signal type_cast_1769_wire : std_logic_vector(15 downto 0);
    signal type_cast_1773_wire : std_logic_vector(15 downto 0);
    signal type_cast_1775_wire : std_logic_vector(15 downto 0);
    signal type_cast_1780_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1788_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1654_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1654_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1654_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1654_resized_base_address <= "00000000000000";
    array_obj_ref_1677_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1677_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1677_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1677_resized_base_address <= "00000000000000";
    ptr_deref_1659_word_offset_0 <= "00000000000000";
    ptr_deref_1681_word_offset_0 <= "00000000000000";
    type_cast_1477_wire_constant <= "00000000000000000000000000010000";
    type_cast_1505_wire_constant <= "1111111111111111";
    type_cast_1516_wire_constant <= "1111111111111111";
    type_cast_1543_wire_constant <= "00000000000000000000000000000010";
    type_cast_1552_wire_constant <= "00000000000000000000000000000000";
    type_cast_1559_wire_constant <= "0000000000000000";
    type_cast_1566_wire_constant <= "0000000000000000";
    type_cast_1573_wire_constant <= "0000000000000000";
    type_cast_1580_wire_constant <= "00000000000000000000000000000100";
    type_cast_1643_wire_constant <= "00000000000000000000000000000010";
    type_cast_1664_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1670_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1691_wire_constant <= "00000000000000000000000000000100";
    type_cast_1709_wire_constant <= "0000000000000100";
    type_cast_1717_wire_constant <= "0000000000000001";
    type_cast_1737_wire_constant <= "0000000000000000";
    type_cast_1763_wire_constant <= "0000000000000000";
    type_cast_1780_wire_constant <= "00000000000000000000000000000001";
    type_cast_1788_wire_constant <= "0000000000000001";
    phi_stmt_1548: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1552_wire_constant & type_cast_1554_wire;
      req <= phi_stmt_1548_req_0 & phi_stmt_1548_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1548",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1548_ack_0,
          idata => idata,
          odata => indvar_1548,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1548
    phi_stmt_1555: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1559_wire_constant & type_cast_1561_wire;
      req <= phi_stmt_1555_req_0 & phi_stmt_1555_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1555",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1555_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1555,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1555
    phi_stmt_1562: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1566_wire_constant & type_cast_1568_wire;
      req <= phi_stmt_1562_req_0 & phi_stmt_1562_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1562",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1562_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1562,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1562
    phi_stmt_1569: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1573_wire_constant & type_cast_1575_wire;
      req <= phi_stmt_1569_req_0 & phi_stmt_1569_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1569",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1569_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1569,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1569
    phi_stmt_1757: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1760_wire & type_cast_1763_wire_constant;
      req <= phi_stmt_1757_req_0 & phi_stmt_1757_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1757",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1757_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1757,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1757
    phi_stmt_1764: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1767_wire & type_cast_1769_wire;
      req <= phi_stmt_1764_req_0 & phi_stmt_1764_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1764",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1764_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1764,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1764
    phi_stmt_1770: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1773_wire & type_cast_1775_wire;
      req <= phi_stmt_1770_req_0 & phi_stmt_1770_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1770",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1770_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1770,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1770
    -- flow-through select operator MUX_1739_inst
    input_dim1x_x2_1740 <= type_cast_1737_wire_constant when (cmp101_1724(0) /=  '0') else inc_1719;
    addr_of_1655_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1655_final_reg_req_0;
      addr_of_1655_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1655_final_reg_req_1;
      addr_of_1655_final_reg_ack_1<= rack(0);
      addr_of_1655_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1655_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1654_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1656,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1678_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1678_final_reg_req_0;
      addr_of_1678_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1678_final_reg_req_1;
      addr_of_1678_final_reg_ack_1<= rack(0);
      addr_of_1678_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1678_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1677_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1679,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1472_inst_req_0;
      type_cast_1472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1472_inst_req_1;
      type_cast_1472_inst_ack_1<= rack(0);
      type_cast_1472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1469,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1485_inst_req_0;
      type_cast_1485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1485_inst_req_1;
      type_cast_1485_inst_ack_1<= rack(0);
      type_cast_1485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1526_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1526_inst_req_0;
      type_cast_1526_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1526_inst_req_1;
      type_cast_1526_inst_ack_1<= rack(0);
      type_cast_1526_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1526_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1527,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1530_inst_req_0;
      type_cast_1530_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1530_inst_req_1;
      type_cast_1530_inst_ack_1<= rack(0);
      type_cast_1530_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1530_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1531,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1534_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1534_inst_req_0;
      type_cast_1534_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1534_inst_req_1;
      type_cast_1534_inst_ack_1<= rack(0);
      type_cast_1534_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1534_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1448,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1535,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1538_inst_req_0;
      type_cast_1538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1538_inst_req_1;
      type_cast_1538_inst_ack_1<= rack(0);
      type_cast_1538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1442,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1554_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1554_inst_req_0;
      type_cast_1554_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1554_inst_req_1;
      type_cast_1554_inst_ack_1<= rack(0);
      type_cast_1554_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1554_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1782,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1554_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1561_inst_req_0;
      type_cast_1561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1561_inst_req_1;
      type_cast_1561_inst_ack_1<= rack(0);
      type_cast_1561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1757,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1561_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1568_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1568_inst_req_0;
      type_cast_1568_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1568_inst_req_1;
      type_cast_1568_inst_ack_1<= rack(0);
      type_cast_1568_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1568_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1568_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1575_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1575_inst_req_0;
      type_cast_1575_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1575_inst_req_1;
      type_cast_1575_inst_ack_1<= rack(0);
      type_cast_1575_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1575_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1770,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1575_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1610_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1610_inst_req_0;
      type_cast_1610_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1610_inst_req_1;
      type_cast_1610_inst_ack_1<= rack(0);
      type_cast_1610_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1610_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1555,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1611,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1614_inst_req_0;
      type_cast_1614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1614_inst_req_1;
      type_cast_1614_inst_ack_1<= rack(0);
      type_cast_1614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1618_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1618_inst_req_0;
      type_cast_1618_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1618_inst_req_1;
      type_cast_1618_inst_ack_1<= rack(0);
      type_cast_1618_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1618_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1597,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1619,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1648_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1648_inst_req_0;
      type_cast_1648_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1648_inst_req_1;
      type_cast_1648_inst_ack_1<= rack(0);
      type_cast_1648_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1648_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1645,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1649,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1686_inst_req_0;
      type_cast_1686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1686_inst_req_1;
      type_cast_1686_inst_ack_1<= rack(0);
      type_cast_1686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1555,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1727_inst_req_0;
      type_cast_1727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1727_inst_req_1;
      type_cast_1727_inst_ack_1<= rack(0);
      type_cast_1727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp101_1724,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc105_1728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1743_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1743_inst_req_0;
      type_cast_1743_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1743_inst_req_1;
      type_cast_1743_inst_ack_1<= rack(0);
      type_cast_1743_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1743_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1733,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1744,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1760_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1760_inst_req_0;
      type_cast_1760_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1760_inst_req_1;
      type_cast_1760_inst_ack_1<= rack(0);
      type_cast_1760_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1760_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add93_1711,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1760_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1767_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1767_inst_req_0;
      type_cast_1767_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1767_inst_req_1;
      type_cast_1767_inst_ack_1<= rack(0);
      type_cast_1767_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1767_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1740,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1767_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1769_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1769_inst_req_0;
      type_cast_1769_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1769_inst_req_1;
      type_cast_1769_inst_ack_1<= rack(0);
      type_cast_1769_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1769_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1562,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1769_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1773_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1773_inst_req_0;
      type_cast_1773_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1773_inst_req_1;
      type_cast_1773_inst_ack_1<= rack(0);
      type_cast_1773_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1773_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1733,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1773_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1775_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1775_inst_req_0;
      type_cast_1775_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1775_inst_req_1;
      type_cast_1775_inst_ack_1<= rack(0);
      type_cast_1775_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1775_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1569,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1775_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1654_index_1_rename
    process(R_idxprom_1653_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1653_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1653_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1654_index_1_resize
    process(idxprom_1649) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1649;
      ov := iv(13 downto 0);
      R_idxprom_1653_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1654_root_address_inst
    process(array_obj_ref_1654_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1654_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1654_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1677_index_1_rename
    process(R_idxprom81_1676_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom81_1676_resized;
      ov(13 downto 0) := iv;
      R_idxprom81_1676_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1677_index_1_resize
    process(idxprom81_1672) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom81_1672;
      ov := iv(13 downto 0);
      R_idxprom81_1676_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1677_root_address_inst
    process(array_obj_ref_1677_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1677_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1677_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1659_addr_0
    process(ptr_deref_1659_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1659_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1659_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1659_base_resize
    process(arrayidx77_1656) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1656;
      ov := iv(13 downto 0);
      ptr_deref_1659_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1659_gather_scatter
    process(ptr_deref_1659_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1659_data_0;
      ov(63 downto 0) := iv;
      tmp78_1660 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1659_root_address_inst
    process(ptr_deref_1659_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1659_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1659_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1681_addr_0
    process(ptr_deref_1681_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1681_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1681_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1681_base_resize
    process(arrayidx82_1679) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1679;
      ov := iv(13 downto 0);
      ptr_deref_1681_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1681_gather_scatter
    process(tmp78_1660) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1660;
      ov(63 downto 0) := iv;
      ptr_deref_1681_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1681_root_address_inst
    process(ptr_deref_1681_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1681_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1681_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1699_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1698;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1699_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1699_branch_req_0,
          ack0 => if_stmt_1699_branch_ack_0,
          ack1 => if_stmt_1699_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1750_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp112_1749;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1750_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1750_branch_req_0,
          ack0 => if_stmt_1750_branch_ack_0,
          ack1 => if_stmt_1750_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1506_inst
    process(call7_1454) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1454, type_cast_1505_wire_constant, tmp_var);
      add41_1507 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1517_inst
    process(call9_1457) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1457, type_cast_1516_wire_constant, tmp_var);
      add54_1518 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1596_inst
    process(sub_1512, mul_1592) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1512, mul_1592, tmp_var);
      sub44_1597 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1606_inst
    process(sub57_1523, mul50_1602) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1523, mul50_1602, tmp_var);
      sub58_1607 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1710_inst
    process(input_dim2x_x1_1555) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1555, type_cast_1709_wire_constant, tmp_var);
      add93_1711 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1718_inst
    process(input_dim1x_x1_1562) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1562, type_cast_1717_wire_constant, tmp_var);
      inc_1719 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1732_inst
    process(inc105_1728, input_dim0x_x2_1569) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc105_1728, input_dim0x_x2_1569, tmp_var);
      inc105x_xinput_dim0x_x2_1733 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1586_inst
    process(add_1491, tmp1_1582) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1491, tmp1_1582, tmp_var);
      add_src_0x_x0_1587 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1692_inst
    process(conv85_1687) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_1687, type_cast_1691_wire_constant, tmp_var);
      add86_1693 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1781_inst
    process(indvar_1548) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1548, type_cast_1780_wire_constant, tmp_var);
      indvarx_xnext_1782 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1628_inst
    process(mul72_1624, conv66_1615) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1624, conv66_1615, tmp_var);
      add73_1629 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1638_inst
    process(mul74_1634, conv61_1611) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1634, conv61_1611, tmp_var);
      add75_1639 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1671_inst
    process(shr80_1666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr80_1666, type_cast_1670_wire_constant, tmp_var);
      idxprom81_1672 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1723_inst
    process(inc_1719, call1_1445) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1719, call1_1445, tmp_var);
      cmp101_1724 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1748_inst
    process(conv107_1744, shr111126_1545) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv107_1744, shr111126_1545, tmp_var);
      cmp112_1749 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1544_inst
    process(conv110_1539) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv110_1539, type_cast_1543_wire_constant, tmp_var);
      shr111126_1545 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1644_inst
    process(add_src_0x_x0_1587) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1587, type_cast_1643_wire_constant, tmp_var);
      shr_1645 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1665_inst
    process(add75_1639) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1639, type_cast_1664_wire_constant, tmp_var);
      shr80_1666 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1591_inst
    process(input_dim0x_x2_1569, call13_1463) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1569, call13_1463, tmp_var);
      mul_1592 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1601_inst
    process(input_dim1x_x1_1562, call13_1463) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1562, call13_1463, tmp_var);
      mul50_1602 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1581_inst
    process(indvar_1548) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1548, type_cast_1580_wire_constant, tmp_var);
      tmp1_1582 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1623_inst
    process(conv71_1619, conv69_1531) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1619, conv69_1531, tmp_var);
      mul72_1624 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1633_inst
    process(add73_1629, conv64_1527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1629, conv64_1527, tmp_var);
      mul74_1634 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1490_inst
    process(shl_1479, conv17_1486) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1479, conv17_1486, tmp_var);
      add_1491 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1478_inst
    process(conv_1473) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1473, type_cast_1477_wire_constant, tmp_var);
      shl_1479 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1511_inst
    process(add41_1507, call14_1466) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1507, call14_1466, tmp_var);
      sub_1512 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1522_inst
    process(add54_1518, call14_1466) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1518, call14_1466, tmp_var);
      sub57_1523 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1697_inst
    process(add86_1693, conv89_1535) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add86_1693, conv89_1535, tmp_var);
      cmp_1698 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1654_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1653_scaled;
      array_obj_ref_1654_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1654_index_offset_req_0;
      array_obj_ref_1654_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1654_index_offset_req_1;
      array_obj_ref_1654_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1677_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom81_1676_scaled;
      array_obj_ref_1677_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1677_index_offset_req_0;
      array_obj_ref_1677_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1677_index_offset_req_1;
      array_obj_ref_1677_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1659_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1659_load_0_req_0;
      ptr_deref_1659_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1659_load_0_req_1;
      ptr_deref_1659_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1659_word_address_0;
      ptr_deref_1659_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1681_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1681_store_0_req_0;
      ptr_deref_1681_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1681_store_0_req_1;
      ptr_deref_1681_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1681_word_address_0;
      data_in <= ptr_deref_1681_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1493_inst RPIPE_Block0_start_1481_inst RPIPE_Block0_start_1496_inst RPIPE_Block0_start_1468_inst RPIPE_Block0_start_1465_inst RPIPE_Block0_start_1462_inst RPIPE_Block0_start_1459_inst RPIPE_Block0_start_1456_inst RPIPE_Block0_start_1453_inst RPIPE_Block0_start_1450_inst RPIPE_Block0_start_1447_inst RPIPE_Block0_start_1444_inst RPIPE_Block0_start_1441_inst RPIPE_Block0_start_1499_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1493_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1481_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1496_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1468_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1465_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1462_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1459_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1456_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1453_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1450_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1447_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1444_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1441_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1499_inst_req_0;
      RPIPE_Block0_start_1493_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1481_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1496_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1468_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1465_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1462_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1459_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1456_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1453_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1450_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1447_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1444_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1441_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1499_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1493_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1481_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1496_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1468_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1465_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1462_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1459_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1456_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1453_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1450_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1447_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1444_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1441_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1499_inst_req_1;
      RPIPE_Block0_start_1493_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1481_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1496_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1468_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1465_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1462_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1459_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1456_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1453_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1450_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1447_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1444_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1441_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1499_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call18_1494 <= data_out(223 downto 208);
      call16_1482 <= data_out(207 downto 192);
      call20_1497 <= data_out(191 downto 176);
      call15_1469 <= data_out(175 downto 160);
      call14_1466 <= data_out(159 downto 144);
      call13_1463 <= data_out(143 downto 128);
      call11_1460 <= data_out(127 downto 112);
      call9_1457 <= data_out(111 downto 96);
      call7_1454 <= data_out(95 downto 80);
      call5_1451 <= data_out(79 downto 64);
      call3_1448 <= data_out(63 downto 48);
      call1_1445 <= data_out(47 downto 32);
      call_1442 <= data_out(31 downto 16);
      call22_1500 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1786_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1786_inst_req_0;
      WPIPE_Block0_done_1786_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1786_inst_req_1;
      WPIPE_Block0_done_1786_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1788_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4641_start: Boolean;
  signal convTransposeB_CP_4641_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1824_inst_ack_0 : boolean;
  signal type_cast_1971_inst_ack_0 : boolean;
  signal type_cast_1828_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1821_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1837_inst_req_1 : boolean;
  signal type_cast_1900_inst_ack_0 : boolean;
  signal type_cast_1841_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1815_inst_ack_1 : boolean;
  signal type_cast_1971_inst_req_0 : boolean;
  signal type_cast_1975_inst_req_1 : boolean;
  signal type_cast_1841_inst_req_0 : boolean;
  signal type_cast_1896_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1824_inst_req_1 : boolean;
  signal type_cast_1828_inst_req_1 : boolean;
  signal type_cast_1888_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1818_inst_req_0 : boolean;
  signal type_cast_1888_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1818_inst_req_1 : boolean;
  signal type_cast_1979_inst_req_1 : boolean;
  signal type_cast_1888_inst_req_1 : boolean;
  signal type_cast_1888_inst_ack_1 : boolean;
  signal type_cast_1828_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1818_inst_ack_1 : boolean;
  signal type_cast_1892_inst_ack_1 : boolean;
  signal type_cast_1975_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1821_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1837_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1849_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1824_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1852_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1837_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1837_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1852_inst_ack_0 : boolean;
  signal type_cast_1896_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1849_inst_req_1 : boolean;
  signal type_cast_2009_inst_req_0 : boolean;
  signal type_cast_1971_inst_req_1 : boolean;
  signal type_cast_1841_inst_req_1 : boolean;
  signal type_cast_1892_inst_req_0 : boolean;
  signal type_cast_1841_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1815_inst_req_1 : boolean;
  signal type_cast_1971_inst_ack_1 : boolean;
  signal array_obj_ref_2015_index_offset_ack_1 : boolean;
  signal type_cast_1892_inst_ack_0 : boolean;
  signal type_cast_1900_inst_req_1 : boolean;
  signal type_cast_1828_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1821_inst_req_1 : boolean;
  signal type_cast_2009_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1815_inst_ack_0 : boolean;
  signal type_cast_1900_inst_ack_1 : boolean;
  signal array_obj_ref_2015_index_offset_ack_0 : boolean;
  signal RPIPE_Block1_start_1818_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1855_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1815_inst_req_0 : boolean;
  signal type_cast_1979_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1855_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1852_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1855_inst_ack_0 : boolean;
  signal type_cast_1896_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1821_inst_ack_1 : boolean;
  signal type_cast_1896_inst_ack_0 : boolean;
  signal type_cast_2009_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1824_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1852_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1855_inst_ack_1 : boolean;
  signal type_cast_1979_inst_req_0 : boolean;
  signal type_cast_1900_inst_req_0 : boolean;
  signal type_cast_1979_inst_ack_0 : boolean;
  signal type_cast_1892_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1849_inst_ack_0 : boolean;
  signal type_cast_1975_inst_ack_0 : boolean;
  signal addr_of_2016_final_reg_req_0 : boolean;
  signal RPIPE_Block1_start_1849_inst_req_0 : boolean;
  signal type_cast_1975_inst_req_0 : boolean;
  signal addr_of_2016_final_reg_req_1 : boolean;
  signal addr_of_2016_final_reg_ack_1 : boolean;
  signal addr_of_2016_final_reg_ack_0 : boolean;
  signal array_obj_ref_2015_index_offset_req_0 : boolean;
  signal array_obj_ref_2015_index_offset_req_1 : boolean;
  signal type_cast_2009_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1797_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1797_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1797_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1797_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1800_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1800_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1800_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1800_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1803_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1803_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1803_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1803_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1806_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1806_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1806_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1806_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1809_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1809_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1809_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1809_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1812_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1812_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1812_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1812_inst_ack_1 : boolean;
  signal ptr_deref_2020_load_0_req_0 : boolean;
  signal ptr_deref_2020_load_0_ack_0 : boolean;
  signal ptr_deref_2020_load_0_req_1 : boolean;
  signal ptr_deref_2020_load_0_ack_1 : boolean;
  signal array_obj_ref_2038_index_offset_req_0 : boolean;
  signal array_obj_ref_2038_index_offset_ack_0 : boolean;
  signal array_obj_ref_2038_index_offset_req_1 : boolean;
  signal array_obj_ref_2038_index_offset_ack_1 : boolean;
  signal addr_of_2039_final_reg_req_0 : boolean;
  signal addr_of_2039_final_reg_ack_0 : boolean;
  signal addr_of_2039_final_reg_req_1 : boolean;
  signal addr_of_2039_final_reg_ack_1 : boolean;
  signal ptr_deref_2042_store_0_req_0 : boolean;
  signal ptr_deref_2042_store_0_ack_0 : boolean;
  signal ptr_deref_2042_store_0_req_1 : boolean;
  signal ptr_deref_2042_store_0_ack_1 : boolean;
  signal type_cast_2047_inst_req_0 : boolean;
  signal type_cast_2047_inst_ack_0 : boolean;
  signal type_cast_2047_inst_req_1 : boolean;
  signal type_cast_2047_inst_ack_1 : boolean;
  signal if_stmt_2060_branch_req_0 : boolean;
  signal if_stmt_2060_branch_ack_1 : boolean;
  signal if_stmt_2060_branch_ack_0 : boolean;
  signal type_cast_2088_inst_req_0 : boolean;
  signal type_cast_2088_inst_ack_0 : boolean;
  signal type_cast_2088_inst_req_1 : boolean;
  signal type_cast_2088_inst_ack_1 : boolean;
  signal type_cast_2104_inst_req_0 : boolean;
  signal type_cast_2104_inst_ack_0 : boolean;
  signal type_cast_2104_inst_req_1 : boolean;
  signal type_cast_2104_inst_ack_1 : boolean;
  signal if_stmt_2111_branch_req_0 : boolean;
  signal if_stmt_2111_branch_ack_1 : boolean;
  signal if_stmt_2111_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2147_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2147_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2147_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2147_inst_ack_1 : boolean;
  signal type_cast_1934_inst_req_0 : boolean;
  signal type_cast_1934_inst_ack_0 : boolean;
  signal type_cast_1934_inst_req_1 : boolean;
  signal type_cast_1934_inst_ack_1 : boolean;
  signal phi_stmt_1931_req_0 : boolean;
  signal phi_stmt_1924_req_0 : boolean;
  signal phi_stmt_1917_req_0 : boolean;
  signal phi_stmt_1910_req_0 : boolean;
  signal type_cast_1936_inst_req_0 : boolean;
  signal type_cast_1936_inst_ack_0 : boolean;
  signal type_cast_1936_inst_req_1 : boolean;
  signal type_cast_1936_inst_ack_1 : boolean;
  signal phi_stmt_1931_req_1 : boolean;
  signal type_cast_1930_inst_req_0 : boolean;
  signal type_cast_1930_inst_ack_0 : boolean;
  signal type_cast_1930_inst_req_1 : boolean;
  signal type_cast_1930_inst_ack_1 : boolean;
  signal phi_stmt_1924_req_1 : boolean;
  signal type_cast_1923_inst_req_0 : boolean;
  signal type_cast_1923_inst_ack_0 : boolean;
  signal type_cast_1923_inst_req_1 : boolean;
  signal type_cast_1923_inst_ack_1 : boolean;
  signal phi_stmt_1917_req_1 : boolean;
  signal type_cast_1916_inst_req_0 : boolean;
  signal type_cast_1916_inst_ack_0 : boolean;
  signal type_cast_1916_inst_req_1 : boolean;
  signal type_cast_1916_inst_ack_1 : boolean;
  signal phi_stmt_1910_req_1 : boolean;
  signal phi_stmt_1910_ack_0 : boolean;
  signal phi_stmt_1917_ack_0 : boolean;
  signal phi_stmt_1924_ack_0 : boolean;
  signal phi_stmt_1931_ack_0 : boolean;
  signal phi_stmt_2118_req_1 : boolean;
  signal type_cast_2134_inst_req_0 : boolean;
  signal type_cast_2134_inst_ack_0 : boolean;
  signal type_cast_2134_inst_req_1 : boolean;
  signal type_cast_2134_inst_ack_1 : boolean;
  signal phi_stmt_2131_req_0 : boolean;
  signal type_cast_2128_inst_req_0 : boolean;
  signal type_cast_2128_inst_ack_0 : boolean;
  signal type_cast_2128_inst_req_1 : boolean;
  signal type_cast_2128_inst_ack_1 : boolean;
  signal phi_stmt_2125_req_0 : boolean;
  signal type_cast_2121_inst_req_0 : boolean;
  signal type_cast_2121_inst_ack_0 : boolean;
  signal type_cast_2121_inst_req_1 : boolean;
  signal type_cast_2121_inst_ack_1 : boolean;
  signal phi_stmt_2118_req_0 : boolean;
  signal type_cast_2136_inst_req_0 : boolean;
  signal type_cast_2136_inst_ack_0 : boolean;
  signal type_cast_2136_inst_req_1 : boolean;
  signal type_cast_2136_inst_ack_1 : boolean;
  signal phi_stmt_2131_req_1 : boolean;
  signal type_cast_2130_inst_req_0 : boolean;
  signal type_cast_2130_inst_ack_0 : boolean;
  signal type_cast_2130_inst_req_1 : boolean;
  signal type_cast_2130_inst_ack_1 : boolean;
  signal phi_stmt_2125_req_1 : boolean;
  signal phi_stmt_2118_ack_0 : boolean;
  signal phi_stmt_2125_ack_0 : boolean;
  signal phi_stmt_2131_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4641_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4641_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4641_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4641_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4641: Block -- control-path 
    signal convTransposeB_CP_4641_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4641_elements(0) <= convTransposeB_CP_4641_start;
    convTransposeB_CP_4641_symbol <= convTransposeB_CP_4641_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1795/$entry
      -- CP-element group 0: 	 branch_block_stmt_1795/branch_block_stmt_1795__entry__
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856__entry__
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/$entry
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_Sample/rr
      -- 
    cr_4834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(0), ack => type_cast_1828_inst_req_1); -- 
    cr_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(0), ack => type_cast_1841_inst_req_1); -- 
    rr_4689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(0), ack => RPIPE_Block1_start_1797_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1795/merge_stmt_2117__exit__
      -- CP-element group 1: 	 branch_block_stmt_1795/assign_stmt_2143__entry__
      -- CP-element group 1: 	 branch_block_stmt_1795/assign_stmt_2143__exit__
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1795/assign_stmt_2143/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/assign_stmt_2143/$exit
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/SplitProtocol/Update/cr
      -- 
    rr_5390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(1), ack => type_cast_1936_inst_req_0); -- 
    cr_5395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(1), ack => type_cast_1936_inst_req_1); -- 
    rr_5413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(1), ack => type_cast_1930_inst_req_0); -- 
    cr_5418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(1), ack => type_cast_1930_inst_req_1); -- 
    rr_5436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(1), ack => type_cast_1923_inst_req_0); -- 
    cr_5441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(1), ack => type_cast_1923_inst_req_1); -- 
    rr_5459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(1), ack => type_cast_1916_inst_req_0); -- 
    cr_5464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(1), ack => type_cast_1916_inst_req_1); -- 
    convTransposeB_CP_4641_elements(1) <= convTransposeB_CP_4641_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_Update/cr
      -- 
    ra_4690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1797_inst_ack_0, ack => convTransposeB_CP_4641_elements(2)); -- 
    cr_4694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(2), ack => RPIPE_Block1_start_1797_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1797_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_Sample/rr
      -- 
    ca_4695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1797_inst_ack_1, ack => convTransposeB_CP_4641_elements(3)); -- 
    rr_4703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(3), ack => RPIPE_Block1_start_1800_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_Update/cr
      -- 
    ra_4704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1800_inst_ack_0, ack => convTransposeB_CP_4641_elements(4)); -- 
    cr_4708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(4), ack => RPIPE_Block1_start_1800_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1800_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_Sample/rr
      -- 
    ca_4709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1800_inst_ack_1, ack => convTransposeB_CP_4641_elements(5)); -- 
    rr_4717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(5), ack => RPIPE_Block1_start_1803_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_Update/cr
      -- 
    ra_4718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1803_inst_ack_0, ack => convTransposeB_CP_4641_elements(6)); -- 
    cr_4722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(6), ack => RPIPE_Block1_start_1803_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1803_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_Sample/rr
      -- 
    ca_4723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1803_inst_ack_1, ack => convTransposeB_CP_4641_elements(7)); -- 
    rr_4731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(7), ack => RPIPE_Block1_start_1806_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_Update/cr
      -- 
    ra_4732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1806_inst_ack_0, ack => convTransposeB_CP_4641_elements(8)); -- 
    cr_4736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(8), ack => RPIPE_Block1_start_1806_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1806_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_Sample/rr
      -- 
    ca_4737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1806_inst_ack_1, ack => convTransposeB_CP_4641_elements(9)); -- 
    rr_4745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(9), ack => RPIPE_Block1_start_1809_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_Update/cr
      -- 
    ra_4746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1809_inst_ack_0, ack => convTransposeB_CP_4641_elements(10)); -- 
    cr_4750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(10), ack => RPIPE_Block1_start_1809_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1809_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_Sample/rr
      -- 
    ca_4751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1809_inst_ack_1, ack => convTransposeB_CP_4641_elements(11)); -- 
    rr_4759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(11), ack => RPIPE_Block1_start_1812_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_Update/cr
      -- 
    ra_4760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1812_inst_ack_0, ack => convTransposeB_CP_4641_elements(12)); -- 
    cr_4764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(12), ack => RPIPE_Block1_start_1812_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1812_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_sample_start_
      -- 
    ca_4765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1812_inst_ack_1, ack => convTransposeB_CP_4641_elements(13)); -- 
    rr_4773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(13), ack => RPIPE_Block1_start_1815_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_update_start_
      -- 
    ra_4774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1815_inst_ack_0, ack => convTransposeB_CP_4641_elements(14)); -- 
    cr_4778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(14), ack => RPIPE_Block1_start_1815_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1815_update_completed_
      -- 
    ca_4779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1815_inst_ack_1, ack => convTransposeB_CP_4641_elements(15)); -- 
    rr_4787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(15), ack => RPIPE_Block1_start_1818_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_sample_completed_
      -- 
    ra_4788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1818_inst_ack_0, ack => convTransposeB_CP_4641_elements(16)); -- 
    cr_4792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(16), ack => RPIPE_Block1_start_1818_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1818_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_sample_start_
      -- 
    ca_4793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1818_inst_ack_1, ack => convTransposeB_CP_4641_elements(17)); -- 
    rr_4801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(17), ack => RPIPE_Block1_start_1821_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_sample_completed_
      -- 
    ra_4802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1821_inst_ack_0, ack => convTransposeB_CP_4641_elements(18)); -- 
    cr_4806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(18), ack => RPIPE_Block1_start_1821_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1821_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_Sample/$entry
      -- 
    ca_4807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1821_inst_ack_1, ack => convTransposeB_CP_4641_elements(19)); -- 
    rr_4815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(19), ack => RPIPE_Block1_start_1824_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_update_start_
      -- 
    ra_4816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1824_inst_ack_0, ack => convTransposeB_CP_4641_elements(20)); -- 
    cr_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(20), ack => RPIPE_Block1_start_1824_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1824_update_completed_
      -- 
    ca_4821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1824_inst_ack_1, ack => convTransposeB_CP_4641_elements(21)); -- 
    rr_4829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(21), ack => type_cast_1828_inst_req_0); -- 
    rr_4843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(21), ack => RPIPE_Block1_start_1837_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_sample_completed_
      -- 
    ra_4830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1828_inst_ack_0, ack => convTransposeB_CP_4641_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1828_update_completed_
      -- 
    ca_4835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1828_inst_ack_1, ack => convTransposeB_CP_4641_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_Update/$entry
      -- 
    ra_4844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1837_inst_ack_0, ack => convTransposeB_CP_4641_elements(24)); -- 
    cr_4848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(24), ack => RPIPE_Block1_start_1837_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1837_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_Sample/$entry
      -- 
    ca_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1837_inst_ack_1, ack => convTransposeB_CP_4641_elements(25)); -- 
    rr_4857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(25), ack => type_cast_1841_inst_req_0); -- 
    rr_4871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(25), ack => RPIPE_Block1_start_1849_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_Sample/$exit
      -- 
    ra_4858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1841_inst_ack_0, ack => convTransposeB_CP_4641_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/type_cast_1841_Update/ca
      -- 
    ca_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1841_inst_ack_1, ack => convTransposeB_CP_4641_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_Sample/$exit
      -- 
    ra_4872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1849_inst_ack_0, ack => convTransposeB_CP_4641_elements(28)); -- 
    cr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(28), ack => RPIPE_Block1_start_1849_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1849_update_completed_
      -- 
    ca_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1849_inst_ack_1, ack => convTransposeB_CP_4641_elements(29)); -- 
    rr_4885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(29), ack => RPIPE_Block1_start_1852_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_Update/cr
      -- 
    ra_4886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1852_inst_ack_0, ack => convTransposeB_CP_4641_elements(30)); -- 
    cr_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(30), ack => RPIPE_Block1_start_1852_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1852_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_sample_start_
      -- 
    ca_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1852_inst_ack_1, ack => convTransposeB_CP_4641_elements(31)); -- 
    rr_4899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(31), ack => RPIPE_Block1_start_1855_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_update_start_
      -- 
    ra_4900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1855_inst_ack_0, ack => convTransposeB_CP_4641_elements(32)); -- 
    cr_4904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(32), ack => RPIPE_Block1_start_1855_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/RPIPE_Block1_start_1855_Update/ca
      -- 
    ca_4905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1855_inst_ack_1, ack => convTransposeB_CP_4641_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/$entry
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856__exit__
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907__entry__
      -- CP-element group 34: 	 branch_block_stmt_1795/assign_stmt_1798_to_assign_stmt_1856/$exit
      -- 
    rr_4944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(34), ack => type_cast_1896_inst_req_0); -- 
    rr_4916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(34), ack => type_cast_1888_inst_req_0); -- 
    cr_4921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(34), ack => type_cast_1888_inst_req_1); -- 
    cr_4949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(34), ack => type_cast_1896_inst_req_1); -- 
    rr_4930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(34), ack => type_cast_1892_inst_req_0); -- 
    cr_4963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(34), ack => type_cast_1900_inst_req_1); -- 
    rr_4958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(34), ack => type_cast_1900_inst_req_0); -- 
    cr_4935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(34), ack => type_cast_1892_inst_req_1); -- 
    convTransposeB_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(23) & convTransposeB_CP_4641_elements(27) & convTransposeB_CP_4641_elements(33);
      gj_convTransposeB_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_Sample/ra
      -- 
    ra_4917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1888_inst_ack_0, ack => convTransposeB_CP_4641_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1888_Update/ca
      -- 
    ca_4922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1888_inst_ack_1, ack => convTransposeB_CP_4641_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_Sample/ra
      -- 
    ra_4931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1892_inst_ack_0, ack => convTransposeB_CP_4641_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1892_Update/$exit
      -- 
    ca_4936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1892_inst_ack_1, ack => convTransposeB_CP_4641_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_sample_completed_
      -- 
    ra_4945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1896_inst_ack_0, ack => convTransposeB_CP_4641_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1896_update_completed_
      -- 
    ca_4950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1896_inst_ack_1, ack => convTransposeB_CP_4641_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_Sample/$exit
      -- 
    ra_4959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1900_inst_ack_0, ack => convTransposeB_CP_4641_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/type_cast_1900_update_completed_
      -- 
    ca_4964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1900_inst_ack_1, ack => convTransposeB_CP_4641_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907/$exit
      -- CP-element group 43: 	 branch_block_stmt_1795/assign_stmt_1863_to_assign_stmt_1907__exit__
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1924/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1917/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1910/$entry
      -- CP-element group 43: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/$entry
      -- 
    rr_5340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(43), ack => type_cast_1934_inst_req_0); -- 
    cr_5345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(43), ack => type_cast_1934_inst_req_1); -- 
    convTransposeB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(36) & convTransposeB_CP_4641_elements(38) & convTransposeB_CP_4641_elements(40) & convTransposeB_CP_4641_elements(42);
      gj_convTransposeB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_sample_completed_
      -- 
    ra_4976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1971_inst_ack_0, ack => convTransposeB_CP_4641_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_update_completed_
      -- 
    ca_4981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1971_inst_ack_1, ack => convTransposeB_CP_4641_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_Sample/$exit
      -- 
    ra_4990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1975_inst_ack_0, ack => convTransposeB_CP_4641_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_update_completed_
      -- 
    ca_4995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1975_inst_ack_1, ack => convTransposeB_CP_4641_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_Sample/ra
      -- 
    ra_5004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1979_inst_ack_0, ack => convTransposeB_CP_4641_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_Update/ca
      -- 
    ca_5009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1979_inst_ack_1, ack => convTransposeB_CP_4641_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_Sample/ra
      -- 
    ra_5018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2009_inst_ack_0, ack => convTransposeB_CP_4641_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_final_index_sum_regn_Sample/req
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_index_resize_1/$entry
      -- 
    ca_5023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2009_inst_ack_1, ack => convTransposeB_CP_4641_elements(51)); -- 
    req_5048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(51), ack => array_obj_ref_2015_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_final_index_sum_regn_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_final_index_sum_regn_Sample/$exit
      -- 
    ack_5049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2015_index_offset_ack_0, ack => convTransposeB_CP_4641_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_request/req
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_root_address_calculated
      -- 
    ack_5054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2015_index_offset_ack_1, ack => convTransposeB_CP_4641_elements(53)); -- 
    req_5063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(53), ack => addr_of_2016_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_request/ack
      -- CP-element group 54: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_sample_completed_
      -- 
    ack_5064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2016_final_reg_ack_0, ack => convTransposeB_CP_4641_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Sample/word_access_start/word_0/rr
      -- 
    ack_5069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2016_final_reg_ack_1, ack => convTransposeB_CP_4641_elements(55)); -- 
    rr_5102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(55), ack => ptr_deref_2020_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Sample/word_access_start/word_0/ra
      -- 
    ra_5103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_load_0_ack_0, ack => convTransposeB_CP_4641_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/ptr_deref_2020_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/ptr_deref_2020_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/ptr_deref_2020_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/ptr_deref_2020_Merge/merge_ack
      -- 
    ca_5114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_load_0_ack_1, ack => convTransposeB_CP_4641_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_final_index_sum_regn_Sample/req
      -- 
    req_5144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(58), ack => array_obj_ref_2038_index_offset_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(45) & convTransposeB_CP_4641_elements(47) & convTransposeB_CP_4641_elements(49);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_final_index_sum_regn_Sample/ack
      -- 
    ack_5145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2038_index_offset_ack_0, ack => convTransposeB_CP_4641_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_request/req
      -- 
    ack_5150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2038_index_offset_ack_1, ack => convTransposeB_CP_4641_elements(60)); -- 
    req_5159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(60), ack => addr_of_2039_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_request/ack
      -- 
    ack_5160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2039_final_reg_ack_0, ack => convTransposeB_CP_4641_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_word_addrgen/root_register_ack
      -- 
    ack_5165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2039_final_reg_ack_1, ack => convTransposeB_CP_4641_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/ptr_deref_2042_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/ptr_deref_2042_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/ptr_deref_2042_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/ptr_deref_2042_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/word_access_start/word_0/rr
      -- 
    rr_5203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(63), ack => ptr_deref_2042_store_0_req_0); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(57) & convTransposeB_CP_4641_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Sample/word_access_start/word_0/ra
      -- 
    ra_5204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_store_0_ack_0, ack => convTransposeB_CP_4641_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Update/word_access_complete/word_0/ca
      -- 
    ca_5215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_store_0_ack_1, ack => convTransposeB_CP_4641_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_Sample/ra
      -- 
    ra_5224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2047_inst_ack_0, ack => convTransposeB_CP_4641_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_Update/ca
      -- 
    ca_5229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2047_inst_ack_1, ack => convTransposeB_CP_4641_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/$exit
      -- CP-element group 68: 	 branch_block_stmt_1795/R_cmp_2061_place
      -- CP-element group 68: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059__exit__
      -- CP-element group 68: 	 branch_block_stmt_1795/if_stmt_2060__entry__
      -- CP-element group 68: 	 branch_block_stmt_1795/if_stmt_2060_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1795/if_stmt_2060_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1795/if_stmt_2060_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1795/if_stmt_2060_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1795/if_stmt_2060_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1795/if_stmt_2060_else_link/$entry
      -- 
    branch_req_5237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(68), ack => if_stmt_2060_branch_req_0); -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(52) & convTransposeB_CP_4641_elements(59) & convTransposeB_CP_4641_elements(65) & convTransposeB_CP_4641_elements(67);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1795/merge_stmt_2066__exit__
      -- CP-element group 69: 	 branch_block_stmt_1795/assign_stmt_2072__entry__
      -- CP-element group 69: 	 branch_block_stmt_1795/assign_stmt_2072__exit__
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128
      -- CP-element group 69: 	 branch_block_stmt_1795/if_stmt_2060_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1795/if_stmt_2060_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1795/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1795/assign_stmt_2072/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/assign_stmt_2072/$exit
      -- CP-element group 69: 	 branch_block_stmt_1795/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1795/merge_stmt_2066_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1795/merge_stmt_2066_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/merge_stmt_2066_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1795/merge_stmt_2066_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2060_branch_ack_1, ack => convTransposeB_CP_4641_elements(69)); -- 
    rr_5574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(69), ack => type_cast_2121_inst_req_0); -- 
    cr_5579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(69), ack => type_cast_2121_inst_req_1); -- 
    rr_5597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(69), ack => type_cast_2136_inst_req_0); -- 
    cr_5602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(69), ack => type_cast_2136_inst_req_1); -- 
    rr_5620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(69), ack => type_cast_2130_inst_req_0); -- 
    cr_5625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(69), ack => type_cast_2130_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1795/merge_stmt_2074__exit__
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110__entry__
      -- CP-element group 70: 	 branch_block_stmt_1795/if_stmt_2060_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1795/if_stmt_2060_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1795/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/$entry
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1795/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1795/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1795/merge_stmt_2074_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1795/merge_stmt_2074_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1795/merge_stmt_2074_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1795/merge_stmt_2074_PhiAck/dummy
      -- 
    else_choice_transition_5246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2060_branch_ack_0, ack => convTransposeB_CP_4641_elements(70)); -- 
    rr_5262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(70), ack => type_cast_2088_inst_req_0); -- 
    cr_5267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(70), ack => type_cast_2088_inst_req_1); -- 
    cr_5281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(70), ack => type_cast_2104_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_Sample/ra
      -- 
    ra_5263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2088_inst_ack_0, ack => convTransposeB_CP_4641_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2088_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_Sample/rr
      -- 
    ca_5268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2088_inst_ack_1, ack => convTransposeB_CP_4641_elements(72)); -- 
    rr_5276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(72), ack => type_cast_2104_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_Sample/ra
      -- 
    ra_5277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2104_inst_ack_0, ack => convTransposeB_CP_4641_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110__exit__
      -- CP-element group 74: 	 branch_block_stmt_1795/if_stmt_2111__entry__
      -- CP-element group 74: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/$exit
      -- CP-element group 74: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1795/assign_stmt_2080_to_assign_stmt_2110/type_cast_2104_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1795/if_stmt_2111_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1795/if_stmt_2111_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1795/if_stmt_2111_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1795/if_stmt_2111_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1795/R_cmp117_2112_place
      -- CP-element group 74: 	 branch_block_stmt_1795/if_stmt_2111_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1795/if_stmt_2111_else_link/$entry
      -- 
    ca_5282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2104_inst_ack_1, ack => convTransposeB_CP_4641_elements(74)); -- 
    branch_req_5290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(74), ack => if_stmt_2111_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1795/merge_stmt_2145__exit__
      -- CP-element group 75: 	 branch_block_stmt_1795/assign_stmt_2150__entry__
      -- CP-element group 75: 	 branch_block_stmt_1795/if_stmt_2111_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1795/if_stmt_2111_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1795/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1795/assign_stmt_2150/$entry
      -- CP-element group 75: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_1795/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1795/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1795/merge_stmt_2145_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1795/merge_stmt_2145_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1795/merge_stmt_2145_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1795/merge_stmt_2145_PhiAck/dummy
      -- 
    if_choice_transition_5295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2111_branch_ack_1, ack => convTransposeB_CP_4641_elements(75)); -- 
    req_5315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(75), ack => WPIPE_Block1_done_2147_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1795/if_stmt_2111_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1795/if_stmt_2111_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2118/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2111_branch_ack_0, ack => convTransposeB_CP_4641_elements(76)); -- 
    rr_5525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(76), ack => type_cast_2134_inst_req_0); -- 
    cr_5530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(76), ack => type_cast_2134_inst_req_1); -- 
    rr_5548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(76), ack => type_cast_2128_inst_req_0); -- 
    cr_5553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(76), ack => type_cast_2128_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_Update/req
      -- 
    ack_5316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2147_inst_ack_0, ack => convTransposeB_CP_4641_elements(77)); -- 
    req_5320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(77), ack => WPIPE_Block1_done_2147_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1795/$exit
      -- CP-element group 78: 	 branch_block_stmt_1795/branch_block_stmt_1795__exit__
      -- CP-element group 78: 	 branch_block_stmt_1795/assign_stmt_2150__exit__
      -- CP-element group 78: 	 branch_block_stmt_1795/return__
      -- CP-element group 78: 	 branch_block_stmt_1795/merge_stmt_2152__exit__
      -- CP-element group 78: 	 branch_block_stmt_1795/assign_stmt_2150/$exit
      -- CP-element group 78: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1795/assign_stmt_2150/WPIPE_Block1_done_2147_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1795/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1795/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1795/merge_stmt_2152_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1795/merge_stmt_2152_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1795/merge_stmt_2152_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1795/merge_stmt_2152_PhiAck/dummy
      -- 
    ack_5321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2147_inst_ack_1, ack => convTransposeB_CP_4641_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/SplitProtocol/Sample/ra
      -- 
    ra_5341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1934_inst_ack_0, ack => convTransposeB_CP_4641_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/SplitProtocol/Update/ca
      -- 
    ca_5346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1934_inst_ack_1, ack => convTransposeB_CP_4641_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/$exit
      -- CP-element group 81: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/$exit
      -- CP-element group 81: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1934/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_req
      -- 
    phi_stmt_1931_req_5347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1931_req_5347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(81), ack => phi_stmt_1931_req_0); -- 
    convTransposeB_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(79) & convTransposeB_CP_4641_elements(80);
      gj_convTransposeB_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1924/$exit
      -- CP-element group 82: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1928_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_req
      -- 
    phi_stmt_1924_req_5355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1924_req_5355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(82), ack => phi_stmt_1924_req_0); -- 
    -- Element group convTransposeB_CP_4641_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeB_CP_4641_elements(43), ack => convTransposeB_CP_4641_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1917/$exit
      -- CP-element group 83: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1921_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_req
      -- 
    phi_stmt_1917_req_5363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1917_req_5363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(83), ack => phi_stmt_1917_req_0); -- 
    -- Element group convTransposeB_CP_4641_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeB_CP_4641_elements(43), ack => convTransposeB_CP_4641_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1910/$exit
      -- CP-element group 84: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1914_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_req
      -- 
    phi_stmt_1910_req_5371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1910_req_5371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(84), ack => phi_stmt_1910_req_0); -- 
    -- Element group convTransposeB_CP_4641_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeB_CP_4641_elements(43), ack => convTransposeB_CP_4641_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1795/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(81) & convTransposeB_CP_4641_elements(82) & convTransposeB_CP_4641_elements(83) & convTransposeB_CP_4641_elements(84);
      gj_convTransposeB_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/SplitProtocol/Sample/ra
      -- 
    ra_5391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1936_inst_ack_0, ack => convTransposeB_CP_4641_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/SplitProtocol/Update/ca
      -- 
    ca_5396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1936_inst_ack_1, ack => convTransposeB_CP_4641_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/$exit
      -- CP-element group 88: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/$exit
      -- CP-element group 88: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_sources/type_cast_1936/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1931/phi_stmt_1931_req
      -- 
    phi_stmt_1931_req_5397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1931_req_5397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(88), ack => phi_stmt_1931_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(86) & convTransposeB_CP_4641_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/SplitProtocol/Sample/ra
      -- 
    ra_5414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1930_inst_ack_0, ack => convTransposeB_CP_4641_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/SplitProtocol/Update/ca
      -- 
    ca_5419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1930_inst_ack_1, ack => convTransposeB_CP_4641_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/$exit
      -- CP-element group 91: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/$exit
      -- CP-element group 91: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_sources/type_cast_1930/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1924/phi_stmt_1924_req
      -- 
    phi_stmt_1924_req_5420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1924_req_5420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(91), ack => phi_stmt_1924_req_1); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(89) & convTransposeB_CP_4641_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/SplitProtocol/Sample/ra
      -- 
    ra_5437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1923_inst_ack_0, ack => convTransposeB_CP_4641_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/SplitProtocol/Update/ca
      -- 
    ca_5442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1923_inst_ack_1, ack => convTransposeB_CP_4641_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/$exit
      -- CP-element group 94: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/$exit
      -- CP-element group 94: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_sources/type_cast_1923/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1917/phi_stmt_1917_req
      -- 
    phi_stmt_1917_req_5443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1917_req_5443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(94), ack => phi_stmt_1917_req_1); -- 
    convTransposeB_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(92) & convTransposeB_CP_4641_elements(93);
      gj_convTransposeB_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/SplitProtocol/Sample/ra
      -- 
    ra_5460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1916_inst_ack_0, ack => convTransposeB_CP_4641_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/SplitProtocol/Update/ca
      -- 
    ca_5465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1916_inst_ack_1, ack => convTransposeB_CP_4641_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/$exit
      -- CP-element group 97: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/$exit
      -- CP-element group 97: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_sources/type_cast_1916/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1910/phi_stmt_1910_req
      -- 
    phi_stmt_1910_req_5466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1910_req_5466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(97), ack => phi_stmt_1910_req_1); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(95) & convTransposeB_CP_4641_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1795/ifx_xend128_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(88) & convTransposeB_CP_4641_elements(91) & convTransposeB_CP_4641_elements(94) & convTransposeB_CP_4641_elements(97);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1795/merge_stmt_1909_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_1795/merge_stmt_1909_PhiAck/$entry
      -- 
    convTransposeB_CP_4641_elements(99) <= OrReduce(convTransposeB_CP_4641_elements(85) & convTransposeB_CP_4641_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1795/merge_stmt_1909_PhiAck/phi_stmt_1910_ack
      -- 
    phi_stmt_1910_ack_5471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1910_ack_0, ack => convTransposeB_CP_4641_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1795/merge_stmt_1909_PhiAck/phi_stmt_1917_ack
      -- 
    phi_stmt_1917_ack_5472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1917_ack_0, ack => convTransposeB_CP_4641_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1795/merge_stmt_1909_PhiAck/phi_stmt_1924_ack
      -- 
    phi_stmt_1924_ack_5473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1924_ack_0, ack => convTransposeB_CP_4641_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1795/merge_stmt_1909_PhiAck/phi_stmt_1931_ack
      -- 
    phi_stmt_1931_ack_5474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1931_ack_0, ack => convTransposeB_CP_4641_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2009_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1979_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2016_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1975_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2015_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1795/merge_stmt_1909__exit__
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059__entry__
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_1971_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2020_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/array_obj_ref_2038_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/addr_of_2039_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/ptr_deref_2042_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1795/assign_stmt_1943_to_assign_stmt_2059/type_cast_2047_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1795/merge_stmt_1909_PhiAck/$exit
      -- 
    rr_4975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => type_cast_1971_inst_req_0); -- 
    cr_4994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => type_cast_1975_inst_req_1); -- 
    cr_5008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => type_cast_1979_inst_req_1); -- 
    rr_5017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => type_cast_2009_inst_req_0); -- 
    cr_4980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => type_cast_1971_inst_req_1); -- 
    cr_5022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => type_cast_2009_inst_req_1); -- 
    rr_5003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => type_cast_1979_inst_req_0); -- 
    rr_4989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => type_cast_1975_inst_req_0); -- 
    req_5068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => addr_of_2016_final_reg_req_1); -- 
    req_5053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => array_obj_ref_2015_index_offset_req_1); -- 
    cr_5113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => ptr_deref_2020_load_0_req_1); -- 
    req_5149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => array_obj_ref_2038_index_offset_req_1); -- 
    req_5164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => addr_of_2039_final_reg_req_1); -- 
    cr_5214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => ptr_deref_2042_store_0_req_1); -- 
    rr_5223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => type_cast_2047_inst_req_0); -- 
    cr_5228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(104), ack => type_cast_2047_inst_req_1); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(100) & convTransposeB_CP_4641_elements(101) & convTransposeB_CP_4641_elements(102) & convTransposeB_CP_4641_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  output  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2118/$exit
      -- CP-element group 105: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2124_konst_delay_trans
      -- CP-element group 105: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_req
      -- 
    phi_stmt_2118_req_5509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2118_req_5509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(105), ack => phi_stmt_2118_req_1); -- 
    -- Element group convTransposeB_CP_4641_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => convTransposeB_CP_4641_elements(76), ack => convTransposeB_CP_4641_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/SplitProtocol/Sample/ra
      -- 
    ra_5526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2134_inst_ack_0, ack => convTransposeB_CP_4641_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/SplitProtocol/Update/ca
      -- 
    ca_5531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2134_inst_ack_1, ack => convTransposeB_CP_4641_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/$exit
      -- CP-element group 108: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/$exit
      -- CP-element group 108: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2134/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_req
      -- 
    phi_stmt_2131_req_5532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2131_req_5532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(108), ack => phi_stmt_2131_req_0); -- 
    convTransposeB_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(106) & convTransposeB_CP_4641_elements(107);
      gj_convTransposeB_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/SplitProtocol/Sample/ra
      -- 
    ra_5549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2128_inst_ack_0, ack => convTransposeB_CP_4641_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/SplitProtocol/Update/ca
      -- 
    ca_5554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2128_inst_ack_1, ack => convTransposeB_CP_4641_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/$exit
      -- CP-element group 111: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/$exit
      -- CP-element group 111: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2128/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_req
      -- 
    phi_stmt_2125_req_5555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2125_req_5555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(111), ack => phi_stmt_2125_req_0); -- 
    convTransposeB_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(109) & convTransposeB_CP_4641_elements(110);
      gj_convTransposeB_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1795/ifx_xelse_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(105) & convTransposeB_CP_4641_elements(108) & convTransposeB_CP_4641_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/SplitProtocol/Sample/ra
      -- 
    ra_5575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2121_inst_ack_0, ack => convTransposeB_CP_4641_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/SplitProtocol/Update/ca
      -- 
    ca_5580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2121_inst_ack_1, ack => convTransposeB_CP_4641_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/$exit
      -- CP-element group 115: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/$exit
      -- CP-element group 115: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_sources/type_cast_2121/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2118/phi_stmt_2118_req
      -- 
    phi_stmt_2118_req_5581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2118_req_5581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(115), ack => phi_stmt_2118_req_0); -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(113) & convTransposeB_CP_4641_elements(114);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/SplitProtocol/Sample/ra
      -- 
    ra_5598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2136_inst_ack_0, ack => convTransposeB_CP_4641_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/SplitProtocol/Update/ca
      -- 
    ca_5603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2136_inst_ack_1, ack => convTransposeB_CP_4641_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/$exit
      -- CP-element group 118: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/$exit
      -- CP-element group 118: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_sources/type_cast_2136/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2131/phi_stmt_2131_req
      -- 
    phi_stmt_2131_req_5604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2131_req_5604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(118), ack => phi_stmt_2131_req_1); -- 
    convTransposeB_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(116) & convTransposeB_CP_4641_elements(117);
      gj_convTransposeB_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/SplitProtocol/Sample/ra
      -- 
    ra_5621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2130_inst_ack_0, ack => convTransposeB_CP_4641_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/SplitProtocol/Update/ca
      -- 
    ca_5626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2130_inst_ack_1, ack => convTransposeB_CP_4641_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/$exit
      -- CP-element group 121: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/$exit
      -- CP-element group 121: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_sources/type_cast_2130/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2125/phi_stmt_2125_req
      -- 
    phi_stmt_2125_req_5627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2125_req_5627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4641_elements(121), ack => phi_stmt_2125_req_1); -- 
    convTransposeB_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(119) & convTransposeB_CP_4641_elements(120);
      gj_convTransposeB_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1795/ifx_xthen_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(115) & convTransposeB_CP_4641_elements(118) & convTransposeB_CP_4641_elements(121);
      gj_convTransposeB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1795/merge_stmt_2117_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_1795/merge_stmt_2117_PhiAck/$entry
      -- 
    convTransposeB_CP_4641_elements(123) <= OrReduce(convTransposeB_CP_4641_elements(112) & convTransposeB_CP_4641_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1795/merge_stmt_2117_PhiAck/phi_stmt_2118_ack
      -- 
    phi_stmt_2118_ack_5632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2118_ack_0, ack => convTransposeB_CP_4641_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1795/merge_stmt_2117_PhiAck/phi_stmt_2125_ack
      -- 
    phi_stmt_2125_ack_5633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2125_ack_0, ack => convTransposeB_CP_4641_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1795/merge_stmt_2117_PhiAck/phi_stmt_2131_ack
      -- 
    phi_stmt_2131_ack_5634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2131_ack_0, ack => convTransposeB_CP_4641_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1795/merge_stmt_2117_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4641_elements(124) & convTransposeB_CP_4641_elements(125) & convTransposeB_CP_4641_elements(126);
      gj_convTransposeB_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4641_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2037_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2037_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2014_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2014_scaled : std_logic_vector(13 downto 0);
    signal add45_1869 : std_logic_vector(15 downto 0);
    signal add58_1880 : std_logic_vector(15 downto 0);
    signal add77_1990 : std_logic_vector(63 downto 0);
    signal add79_2000 : std_logic_vector(63 downto 0);
    signal add91_2054 : std_logic_vector(31 downto 0);
    signal add98_2072 : std_logic_vector(15 downto 0);
    signal add_1847 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1948 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2015_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2015_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2015_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2015_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2015_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2015_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2038_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2038_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2038_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2038_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2038_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2038_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2017 : std_logic_vector(31 downto 0);
    signal arrayidx87_2040 : std_logic_vector(31 downto 0);
    signal call11_1816 : std_logic_vector(15 downto 0);
    signal call13_1819 : std_logic_vector(15 downto 0);
    signal call14_1822 : std_logic_vector(15 downto 0);
    signal call15_1825 : std_logic_vector(15 downto 0);
    signal call16_1838 : std_logic_vector(15 downto 0);
    signal call18_1850 : std_logic_vector(15 downto 0);
    signal call1_1801 : std_logic_vector(15 downto 0);
    signal call20_1853 : std_logic_vector(15 downto 0);
    signal call22_1856 : std_logic_vector(15 downto 0);
    signal call3_1804 : std_logic_vector(15 downto 0);
    signal call5_1807 : std_logic_vector(15 downto 0);
    signal call7_1810 : std_logic_vector(15 downto 0);
    signal call9_1813 : std_logic_vector(15 downto 0);
    signal call_1798 : std_logic_vector(15 downto 0);
    signal cmp106_2085 : std_logic_vector(0 downto 0);
    signal cmp117_2110 : std_logic_vector(0 downto 0);
    signal cmp_2059 : std_logic_vector(0 downto 0);
    signal conv112_2105 : std_logic_vector(31 downto 0);
    signal conv115_1901 : std_logic_vector(31 downto 0);
    signal conv17_1842 : std_logic_vector(31 downto 0);
    signal conv65_1972 : std_logic_vector(63 downto 0);
    signal conv68_1889 : std_logic_vector(63 downto 0);
    signal conv70_1976 : std_logic_vector(63 downto 0);
    signal conv73_1893 : std_logic_vector(63 downto 0);
    signal conv75_1980 : std_logic_vector(63 downto 0);
    signal conv90_2048 : std_logic_vector(31 downto 0);
    signal conv94_1897 : std_logic_vector(31 downto 0);
    signal conv_1829 : std_logic_vector(31 downto 0);
    signal idxprom86_2033 : std_logic_vector(63 downto 0);
    signal idxprom_2010 : std_logic_vector(63 downto 0);
    signal inc110_2089 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2094 : std_logic_vector(15 downto 0);
    signal inc_2080 : std_logic_vector(15 downto 0);
    signal indvar_1910 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2143 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2131 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1931 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2125 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1924 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2101 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2118 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1917 : std_logic_vector(15 downto 0);
    signal mul54_1963 : std_logic_vector(15 downto 0);
    signal mul76_1985 : std_logic_vector(63 downto 0);
    signal mul78_1995 : std_logic_vector(63 downto 0);
    signal mul_1953 : std_logic_vector(15 downto 0);
    signal ptr_deref_2020_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2020_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2042_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2042_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1835 : std_logic_vector(31 downto 0);
    signal shr116132_1907 : std_logic_vector(31 downto 0);
    signal shr131_1863 : std_logic_vector(15 downto 0);
    signal shr81_2006 : std_logic_vector(31 downto 0);
    signal shr85_2027 : std_logic_vector(63 downto 0);
    signal sub48_1958 : std_logic_vector(15 downto 0);
    signal sub61_1885 : std_logic_vector(15 downto 0);
    signal sub62_1968 : std_logic_vector(15 downto 0);
    signal sub_1874 : std_logic_vector(15 downto 0);
    signal tmp1_1943 : std_logic_vector(31 downto 0);
    signal tmp83_2021 : std_logic_vector(63 downto 0);
    signal type_cast_1833_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1861_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1867_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1878_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1905_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1914_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1916_wire : std_logic_vector(31 downto 0);
    signal type_cast_1921_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1923_wire : std_logic_vector(15 downto 0);
    signal type_cast_1928_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1930_wire : std_logic_vector(15 downto 0);
    signal type_cast_1934_wire : std_logic_vector(15 downto 0);
    signal type_cast_1936_wire : std_logic_vector(15 downto 0);
    signal type_cast_1941_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2004_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2025_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2031_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2052_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2070_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2078_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2098_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2121_wire : std_logic_vector(15 downto 0);
    signal type_cast_2124_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2128_wire : std_logic_vector(15 downto 0);
    signal type_cast_2130_wire : std_logic_vector(15 downto 0);
    signal type_cast_2134_wire : std_logic_vector(15 downto 0);
    signal type_cast_2136_wire : std_logic_vector(15 downto 0);
    signal type_cast_2141_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2149_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2015_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2015_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2015_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2015_resized_base_address <= "00000000000000";
    array_obj_ref_2038_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2038_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2038_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2038_resized_base_address <= "00000000000000";
    ptr_deref_2020_word_offset_0 <= "00000000000000";
    ptr_deref_2042_word_offset_0 <= "00000000000000";
    type_cast_1833_wire_constant <= "00000000000000000000000000010000";
    type_cast_1861_wire_constant <= "0000000000000010";
    type_cast_1867_wire_constant <= "1111111111111111";
    type_cast_1878_wire_constant <= "1111111111111111";
    type_cast_1905_wire_constant <= "00000000000000000000000000000001";
    type_cast_1914_wire_constant <= "00000000000000000000000000000000";
    type_cast_1921_wire_constant <= "0000000000000000";
    type_cast_1928_wire_constant <= "0000000000000000";
    type_cast_1941_wire_constant <= "00000000000000000000000000000100";
    type_cast_2004_wire_constant <= "00000000000000000000000000000010";
    type_cast_2025_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2031_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2052_wire_constant <= "00000000000000000000000000000100";
    type_cast_2070_wire_constant <= "0000000000000100";
    type_cast_2078_wire_constant <= "0000000000000001";
    type_cast_2098_wire_constant <= "0000000000000000";
    type_cast_2124_wire_constant <= "0000000000000000";
    type_cast_2141_wire_constant <= "00000000000000000000000000000001";
    type_cast_2149_wire_constant <= "0000000000000001";
    phi_stmt_1910: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1914_wire_constant & type_cast_1916_wire;
      req <= phi_stmt_1910_req_0 & phi_stmt_1910_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1910",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1910_ack_0,
          idata => idata,
          odata => indvar_1910,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1910
    phi_stmt_1917: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1921_wire_constant & type_cast_1923_wire;
      req <= phi_stmt_1917_req_0 & phi_stmt_1917_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1917",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1917_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1917,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1917
    phi_stmt_1924: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1928_wire_constant & type_cast_1930_wire;
      req <= phi_stmt_1924_req_0 & phi_stmt_1924_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1924",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1924_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1924,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1924
    phi_stmt_1931: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1934_wire & type_cast_1936_wire;
      req <= phi_stmt_1931_req_0 & phi_stmt_1931_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1931",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1931_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1931,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1931
    phi_stmt_2118: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2121_wire & type_cast_2124_wire_constant;
      req <= phi_stmt_2118_req_0 & phi_stmt_2118_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2118",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2118_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2118,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2118
    phi_stmt_2125: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2128_wire & type_cast_2130_wire;
      req <= phi_stmt_2125_req_0 & phi_stmt_2125_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2125",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2125_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2125,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2125
    phi_stmt_2131: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2134_wire & type_cast_2136_wire;
      req <= phi_stmt_2131_req_0 & phi_stmt_2131_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2131",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2131_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2131,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2131
    -- flow-through select operator MUX_2100_inst
    input_dim1x_x2_2101 <= type_cast_2098_wire_constant when (cmp106_2085(0) /=  '0') else inc_2080;
    addr_of_2016_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2016_final_reg_req_0;
      addr_of_2016_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2016_final_reg_req_1;
      addr_of_2016_final_reg_ack_1<= rack(0);
      addr_of_2016_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2016_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2015_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2017,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2039_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2039_final_reg_req_0;
      addr_of_2039_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2039_final_reg_req_1;
      addr_of_2039_final_reg_ack_1<= rack(0);
      addr_of_2039_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2039_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2038_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2040,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1828_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1828_inst_req_0;
      type_cast_1828_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1828_inst_req_1;
      type_cast_1828_inst_ack_1<= rack(0);
      type_cast_1828_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1828_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1825,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1829,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1841_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1841_inst_req_0;
      type_cast_1841_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1841_inst_req_1;
      type_cast_1841_inst_ack_1<= rack(0);
      type_cast_1841_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1841_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1838,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1842,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1888_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1888_inst_req_0;
      type_cast_1888_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1888_inst_req_1;
      type_cast_1888_inst_ack_1<= rack(0);
      type_cast_1888_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1888_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1856,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_1889,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1892_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1892_inst_req_0;
      type_cast_1892_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1892_inst_req_1;
      type_cast_1892_inst_ack_1<= rack(0);
      type_cast_1892_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1892_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1853,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1893,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1896_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1896_inst_req_0;
      type_cast_1896_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1896_inst_req_1;
      type_cast_1896_inst_ack_1<= rack(0);
      type_cast_1896_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1896_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1804,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1897,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1900_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1900_inst_req_0;
      type_cast_1900_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1900_inst_req_1;
      type_cast_1900_inst_ack_1<= rack(0);
      type_cast_1900_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1900_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1901,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1916_inst_req_0;
      type_cast_1916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1916_inst_req_1;
      type_cast_1916_inst_ack_1<= rack(0);
      type_cast_1916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1916_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1923_inst_req_0;
      type_cast_1923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1923_inst_req_1;
      type_cast_1923_inst_ack_1<= rack(0);
      type_cast_1923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2118,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1923_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1930_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1930_inst_req_0;
      type_cast_1930_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1930_inst_req_1;
      type_cast_1930_inst_ack_1<= rack(0);
      type_cast_1930_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1930_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1930_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1934_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1934_inst_req_0;
      type_cast_1934_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1934_inst_req_1;
      type_cast_1934_inst_ack_1<= rack(0);
      type_cast_1934_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1934_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr131_1863,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1934_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1936_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1936_inst_req_0;
      type_cast_1936_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1936_inst_req_1;
      type_cast_1936_inst_ack_1<= rack(0);
      type_cast_1936_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1936_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2131,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1936_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1971_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1971_inst_req_0;
      type_cast_1971_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1971_inst_req_1;
      type_cast_1971_inst_ack_1<= rack(0);
      type_cast_1971_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1971_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_1972,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1975_inst_req_0;
      type_cast_1975_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1975_inst_req_1;
      type_cast_1975_inst_ack_1<= rack(0);
      type_cast_1975_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1975_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_1968,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_1976,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1979_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1979_inst_req_0;
      type_cast_1979_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1979_inst_req_1;
      type_cast_1979_inst_ack_1<= rack(0);
      type_cast_1979_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1979_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_1958,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_1980,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2009_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2009_inst_req_0;
      type_cast_2009_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2009_inst_req_1;
      type_cast_2009_inst_ack_1<= rack(0);
      type_cast_2009_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2009_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2010,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2047_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2047_inst_req_0;
      type_cast_2047_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2047_inst_req_1;
      type_cast_2047_inst_ack_1<= rack(0);
      type_cast_2047_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2047_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2048,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2088_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2088_inst_req_0;
      type_cast_2088_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2088_inst_req_1;
      type_cast_2088_inst_ack_1<= rack(0);
      type_cast_2088_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2088_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2085,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2089,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2104_inst_req_0;
      type_cast_2104_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2104_inst_req_1;
      type_cast_2104_inst_ack_1<= rack(0);
      type_cast_2104_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2104_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2094,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2105,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2121_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2121_inst_req_0;
      type_cast_2121_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2121_inst_req_1;
      type_cast_2121_inst_ack_1<= rack(0);
      type_cast_2121_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2121_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2072,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2121_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2128_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2128_inst_req_0;
      type_cast_2128_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2128_inst_req_1;
      type_cast_2128_inst_ack_1<= rack(0);
      type_cast_2128_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2128_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2128_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2130_inst_req_0;
      type_cast_2130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2130_inst_req_1;
      type_cast_2130_inst_ack_1<= rack(0);
      type_cast_2130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2130_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1924,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2130_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2134_inst_req_0;
      type_cast_2134_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2134_inst_req_1;
      type_cast_2134_inst_ack_1<= rack(0);
      type_cast_2134_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2134_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2094,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2134_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2136_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2136_inst_req_0;
      type_cast_2136_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2136_inst_req_1;
      type_cast_2136_inst_ack_1<= rack(0);
      type_cast_2136_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2136_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1931,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2136_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2015_index_1_rename
    process(R_idxprom_2014_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2014_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2014_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2015_index_1_resize
    process(idxprom_2010) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2010;
      ov := iv(13 downto 0);
      R_idxprom_2014_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2015_root_address_inst
    process(array_obj_ref_2015_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2015_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2015_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2038_index_1_rename
    process(R_idxprom86_2037_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2037_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2037_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2038_index_1_resize
    process(idxprom86_2033) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2033;
      ov := iv(13 downto 0);
      R_idxprom86_2037_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2038_root_address_inst
    process(array_obj_ref_2038_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2038_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2038_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2020_addr_0
    process(ptr_deref_2020_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2020_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2020_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2020_base_resize
    process(arrayidx82_2017) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2017;
      ov := iv(13 downto 0);
      ptr_deref_2020_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2020_gather_scatter
    process(ptr_deref_2020_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2020_data_0;
      ov(63 downto 0) := iv;
      tmp83_2021 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2020_root_address_inst
    process(ptr_deref_2020_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2020_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2020_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2042_addr_0
    process(ptr_deref_2042_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2042_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2042_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2042_base_resize
    process(arrayidx87_2040) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2040;
      ov := iv(13 downto 0);
      ptr_deref_2042_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2042_gather_scatter
    process(tmp83_2021) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2021;
      ov(63 downto 0) := iv;
      ptr_deref_2042_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2042_root_address_inst
    process(ptr_deref_2042_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2042_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2042_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2060_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2059;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2060_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2060_branch_req_0,
          ack0 => if_stmt_2060_branch_ack_0,
          ack1 => if_stmt_2060_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2111_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp117_2110;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2111_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2111_branch_req_0,
          ack0 => if_stmt_2111_branch_ack_0,
          ack1 => if_stmt_2111_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1868_inst
    process(call7_1810) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1810, type_cast_1867_wire_constant, tmp_var);
      add45_1869 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1879_inst
    process(call9_1813) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1813, type_cast_1878_wire_constant, tmp_var);
      add58_1880 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1957_inst
    process(sub_1874, mul_1953) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1874, mul_1953, tmp_var);
      sub48_1958 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1967_inst
    process(sub61_1885, mul54_1963) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_1885, mul54_1963, tmp_var);
      sub62_1968 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2071_inst
    process(input_dim2x_x1_1917) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1917, type_cast_2070_wire_constant, tmp_var);
      add98_2072 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2079_inst
    process(input_dim1x_x1_1924) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1924, type_cast_2078_wire_constant, tmp_var);
      inc_2080 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2093_inst
    process(inc110_2089, input_dim0x_x2_1931) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2089, input_dim0x_x2_1931, tmp_var);
      inc110x_xinput_dim0x_x2_2094 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1947_inst
    process(add_1847, tmp1_1943) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1847, tmp1_1943, tmp_var);
      add_src_0x_x0_1948 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2053_inst
    process(conv90_2048) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2048, type_cast_2052_wire_constant, tmp_var);
      add91_2054 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2142_inst
    process(indvar_1910) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1910, type_cast_2141_wire_constant, tmp_var);
      indvarx_xnext_2143 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1989_inst
    process(mul76_1985, conv70_1976) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_1985, conv70_1976, tmp_var);
      add77_1990 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1999_inst
    process(mul78_1995, conv65_1972) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_1995, conv65_1972, tmp_var);
      add79_2000 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2032_inst
    process(shr85_2027) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2027, type_cast_2031_wire_constant, tmp_var);
      idxprom86_2033 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2084_inst
    process(inc_2080, call1_1801) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2080, call1_1801, tmp_var);
      cmp106_2085 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2109_inst
    process(conv112_2105, shr116132_1907) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2105, shr116132_1907, tmp_var);
      cmp117_2110 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1862_inst
    process(call_1798) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1798, type_cast_1861_wire_constant, tmp_var);
      shr131_1863 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1906_inst
    process(conv115_1901) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_1901, type_cast_1905_wire_constant, tmp_var);
      shr116132_1907 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2005_inst
    process(add_src_0x_x0_1948) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1948, type_cast_2004_wire_constant, tmp_var);
      shr81_2006 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2026_inst
    process(add79_2000) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2000, type_cast_2025_wire_constant, tmp_var);
      shr85_2027 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1952_inst
    process(input_dim0x_x2_1931, call13_1819) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1931, call13_1819, tmp_var);
      mul_1953 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1962_inst
    process(input_dim1x_x1_1924, call13_1819) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1924, call13_1819, tmp_var);
      mul54_1963 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1942_inst
    process(indvar_1910) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1910, type_cast_1941_wire_constant, tmp_var);
      tmp1_1943 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1984_inst
    process(conv75_1980, conv73_1893) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_1980, conv73_1893, tmp_var);
      mul76_1985 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1994_inst
    process(add77_1990, conv68_1889) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_1990, conv68_1889, tmp_var);
      mul78_1995 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1846_inst
    process(shl_1835, conv17_1842) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1835, conv17_1842, tmp_var);
      add_1847 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1834_inst
    process(conv_1829) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1829, type_cast_1833_wire_constant, tmp_var);
      shl_1835 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1873_inst
    process(add45_1869, call14_1822) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_1869, call14_1822, tmp_var);
      sub_1874 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1884_inst
    process(add58_1880, call14_1822) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_1880, call14_1822, tmp_var);
      sub61_1885 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2058_inst
    process(add91_2054, conv94_1897) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2054, conv94_1897, tmp_var);
      cmp_2059 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2015_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2014_scaled;
      array_obj_ref_2015_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2015_index_offset_req_0;
      array_obj_ref_2015_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2015_index_offset_req_1;
      array_obj_ref_2015_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2038_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2037_scaled;
      array_obj_ref_2038_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2038_index_offset_req_0;
      array_obj_ref_2038_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2038_index_offset_req_1;
      array_obj_ref_2038_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : ptr_deref_2020_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2020_load_0_req_0;
      ptr_deref_2020_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2020_load_0_req_1;
      ptr_deref_2020_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2020_word_address_0;
      ptr_deref_2020_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2042_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2042_store_0_req_0;
      ptr_deref_2042_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2042_store_0_req_1;
      ptr_deref_2042_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2042_word_address_0;
      data_in <= ptr_deref_2042_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1849_inst RPIPE_Block1_start_1852_inst RPIPE_Block1_start_1855_inst RPIPE_Block1_start_1837_inst RPIPE_Block1_start_1824_inst RPIPE_Block1_start_1821_inst RPIPE_Block1_start_1818_inst RPIPE_Block1_start_1815_inst RPIPE_Block1_start_1812_inst RPIPE_Block1_start_1809_inst RPIPE_Block1_start_1806_inst RPIPE_Block1_start_1803_inst RPIPE_Block1_start_1800_inst RPIPE_Block1_start_1797_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block1_start_1849_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_1852_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1855_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1837_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1824_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1821_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1818_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1815_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1812_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1809_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1806_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1803_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1800_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1797_inst_req_0;
      RPIPE_Block1_start_1849_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_1852_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1855_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1837_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1824_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1821_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1818_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1815_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1812_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1809_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1806_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1803_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1800_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1797_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block1_start_1849_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_1852_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1855_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1837_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1824_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1821_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1818_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1815_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1812_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1809_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1806_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1803_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1800_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1797_inst_req_1;
      RPIPE_Block1_start_1849_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_1852_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1855_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1837_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1824_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1821_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1818_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1815_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1812_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1809_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1806_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1803_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1800_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1797_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call18_1850 <= data_out(223 downto 208);
      call20_1853 <= data_out(207 downto 192);
      call22_1856 <= data_out(191 downto 176);
      call16_1838 <= data_out(175 downto 160);
      call15_1825 <= data_out(159 downto 144);
      call14_1822 <= data_out(143 downto 128);
      call13_1819 <= data_out(127 downto 112);
      call11_1816 <= data_out(111 downto 96);
      call9_1813 <= data_out(95 downto 80);
      call7_1810 <= data_out(79 downto 64);
      call5_1807 <= data_out(63 downto 48);
      call3_1804 <= data_out(47 downto 32);
      call1_1801 <= data_out(31 downto 16);
      call_1798 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2147_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2147_inst_req_0;
      WPIPE_Block1_done_2147_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2147_inst_req_1;
      WPIPE_Block1_done_2147_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2149_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5651_start: Boolean;
  signal convTransposeC_CP_5651_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2261_inst_req_1 : boolean;
  signal type_cast_2249_inst_req_0 : boolean;
  signal type_cast_2202_inst_ack_0 : boolean;
  signal type_cast_2261_inst_ack_0 : boolean;
  signal type_cast_2347_inst_ack_0 : boolean;
  signal type_cast_2343_inst_req_1 : boolean;
  signal array_obj_ref_2410_index_offset_req_0 : boolean;
  signal array_obj_ref_2410_index_offset_ack_0 : boolean;
  signal type_cast_2347_inst_req_1 : boolean;
  signal type_cast_2347_inst_req_0 : boolean;
  signal type_cast_2202_inst_ack_1 : boolean;
  signal type_cast_2249_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2213_inst_req_1 : boolean;
  signal type_cast_2261_inst_ack_1 : boolean;
  signal type_cast_2351_inst_ack_0 : boolean;
  signal type_cast_2253_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2198_inst_req_0 : boolean;
  signal type_cast_2351_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2198_inst_ack_0 : boolean;
  signal type_cast_2381_inst_req_0 : boolean;
  signal type_cast_2381_inst_ack_0 : boolean;
  signal type_cast_2257_inst_req_0 : boolean;
  signal type_cast_2257_inst_ack_0 : boolean;
  signal type_cast_2381_inst_req_1 : boolean;
  signal type_cast_2381_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2213_inst_ack_1 : boolean;
  signal array_obj_ref_2387_index_offset_req_0 : boolean;
  signal type_cast_2257_inst_req_1 : boolean;
  signal type_cast_2343_inst_ack_0 : boolean;
  signal array_obj_ref_2387_index_offset_ack_0 : boolean;
  signal type_cast_2261_inst_req_0 : boolean;
  signal type_cast_2257_inst_ack_1 : boolean;
  signal array_obj_ref_2387_index_offset_req_1 : boolean;
  signal type_cast_2253_inst_ack_1 : boolean;
  signal array_obj_ref_2387_index_offset_ack_1 : boolean;
  signal RPIPE_Block2_start_2198_inst_req_1 : boolean;
  signal type_cast_2202_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2198_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2216_inst_ack_0 : boolean;
  signal type_cast_2343_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2216_inst_req_1 : boolean;
  signal array_obj_ref_2410_index_offset_req_1 : boolean;
  signal array_obj_ref_2410_index_offset_ack_1 : boolean;
  signal type_cast_2253_inst_ack_0 : boolean;
  signal addr_of_2388_final_reg_ack_0 : boolean;
  signal RPIPE_Block2_start_2213_inst_req_0 : boolean;
  signal type_cast_2189_inst_req_1 : boolean;
  signal addr_of_2388_final_reg_ack_1 : boolean;
  signal RPIPE_Block2_start_2216_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2213_inst_ack_0 : boolean;
  signal type_cast_2343_inst_ack_1 : boolean;
  signal ptr_deref_2392_load_0_req_0 : boolean;
  signal ptr_deref_2392_load_0_ack_0 : boolean;
  signal RPIPE_Block2_start_2216_inst_ack_1 : boolean;
  signal type_cast_2189_inst_ack_1 : boolean;
  signal ptr_deref_2392_load_0_req_1 : boolean;
  signal addr_of_2388_final_reg_req_1 : boolean;
  signal type_cast_2253_inst_req_0 : boolean;
  signal addr_of_2411_final_reg_req_1 : boolean;
  signal addr_of_2411_final_reg_ack_1 : boolean;
  signal ptr_deref_2392_load_0_ack_1 : boolean;
  signal type_cast_2351_inst_ack_1 : boolean;
  signal addr_of_2411_final_reg_req_0 : boolean;
  signal addr_of_2411_final_reg_ack_0 : boolean;
  signal addr_of_2388_final_reg_req_0 : boolean;
  signal type_cast_2249_inst_ack_1 : boolean;
  signal type_cast_2351_inst_req_1 : boolean;
  signal type_cast_2202_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2210_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2210_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2210_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2210_inst_req_0 : boolean;
  signal type_cast_2249_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2158_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2158_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2158_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2158_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2161_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2161_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2161_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2161_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2164_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2164_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2164_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2164_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2167_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2167_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2167_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2167_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2170_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2170_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2170_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2170_inst_ack_1 : boolean;
  signal type_cast_2347_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2173_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2173_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2173_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2173_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2176_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2176_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2176_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2176_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2179_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2179_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2179_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2179_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2182_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2182_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2182_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2182_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2185_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2185_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2185_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2185_inst_ack_1 : boolean;
  signal type_cast_2189_inst_req_0 : boolean;
  signal type_cast_2189_inst_ack_0 : boolean;
  signal ptr_deref_2414_store_0_req_0 : boolean;
  signal ptr_deref_2414_store_0_ack_0 : boolean;
  signal ptr_deref_2414_store_0_req_1 : boolean;
  signal ptr_deref_2414_store_0_ack_1 : boolean;
  signal type_cast_2419_inst_req_0 : boolean;
  signal type_cast_2419_inst_ack_0 : boolean;
  signal type_cast_2419_inst_req_1 : boolean;
  signal type_cast_2419_inst_ack_1 : boolean;
  signal if_stmt_2432_branch_req_0 : boolean;
  signal if_stmt_2432_branch_ack_1 : boolean;
  signal if_stmt_2432_branch_ack_0 : boolean;
  signal type_cast_2460_inst_req_0 : boolean;
  signal type_cast_2460_inst_ack_0 : boolean;
  signal type_cast_2460_inst_req_1 : boolean;
  signal type_cast_2460_inst_ack_1 : boolean;
  signal type_cast_2476_inst_req_0 : boolean;
  signal type_cast_2476_inst_ack_0 : boolean;
  signal type_cast_2476_inst_req_1 : boolean;
  signal type_cast_2476_inst_ack_1 : boolean;
  signal if_stmt_2483_branch_req_0 : boolean;
  signal if_stmt_2483_branch_ack_1 : boolean;
  signal if_stmt_2483_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2519_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2519_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2519_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2519_inst_ack_1 : boolean;
  signal phi_stmt_2282_req_0 : boolean;
  signal phi_stmt_2289_req_0 : boolean;
  signal phi_stmt_2296_req_0 : boolean;
  signal type_cast_2306_inst_req_0 : boolean;
  signal type_cast_2306_inst_ack_0 : boolean;
  signal type_cast_2306_inst_req_1 : boolean;
  signal type_cast_2306_inst_ack_1 : boolean;
  signal phi_stmt_2303_req_0 : boolean;
  signal type_cast_2288_inst_req_0 : boolean;
  signal type_cast_2288_inst_ack_0 : boolean;
  signal type_cast_2288_inst_req_1 : boolean;
  signal type_cast_2288_inst_ack_1 : boolean;
  signal phi_stmt_2282_req_1 : boolean;
  signal type_cast_2295_inst_req_0 : boolean;
  signal type_cast_2295_inst_ack_0 : boolean;
  signal type_cast_2295_inst_req_1 : boolean;
  signal type_cast_2295_inst_ack_1 : boolean;
  signal phi_stmt_2289_req_1 : boolean;
  signal type_cast_2302_inst_req_0 : boolean;
  signal type_cast_2302_inst_ack_0 : boolean;
  signal type_cast_2302_inst_req_1 : boolean;
  signal type_cast_2302_inst_ack_1 : boolean;
  signal phi_stmt_2296_req_1 : boolean;
  signal type_cast_2308_inst_req_0 : boolean;
  signal type_cast_2308_inst_ack_0 : boolean;
  signal type_cast_2308_inst_req_1 : boolean;
  signal type_cast_2308_inst_ack_1 : boolean;
  signal phi_stmt_2303_req_1 : boolean;
  signal phi_stmt_2282_ack_0 : boolean;
  signal phi_stmt_2289_ack_0 : boolean;
  signal phi_stmt_2296_ack_0 : boolean;
  signal phi_stmt_2303_ack_0 : boolean;
  signal phi_stmt_2490_req_1 : boolean;
  signal type_cast_2500_inst_req_0 : boolean;
  signal type_cast_2500_inst_ack_0 : boolean;
  signal type_cast_2500_inst_req_1 : boolean;
  signal type_cast_2500_inst_ack_1 : boolean;
  signal phi_stmt_2497_req_0 : boolean;
  signal type_cast_2506_inst_req_0 : boolean;
  signal type_cast_2506_inst_ack_0 : boolean;
  signal type_cast_2506_inst_req_1 : boolean;
  signal type_cast_2506_inst_ack_1 : boolean;
  signal phi_stmt_2503_req_0 : boolean;
  signal type_cast_2493_inst_req_0 : boolean;
  signal type_cast_2493_inst_ack_0 : boolean;
  signal type_cast_2493_inst_req_1 : boolean;
  signal type_cast_2493_inst_ack_1 : boolean;
  signal phi_stmt_2490_req_0 : boolean;
  signal type_cast_2502_inst_req_0 : boolean;
  signal type_cast_2502_inst_ack_0 : boolean;
  signal type_cast_2502_inst_req_1 : boolean;
  signal type_cast_2502_inst_ack_1 : boolean;
  signal phi_stmt_2497_req_1 : boolean;
  signal type_cast_2508_inst_req_0 : boolean;
  signal type_cast_2508_inst_ack_0 : boolean;
  signal type_cast_2508_inst_req_1 : boolean;
  signal type_cast_2508_inst_ack_1 : boolean;
  signal phi_stmt_2503_req_1 : boolean;
  signal phi_stmt_2490_ack_0 : boolean;
  signal phi_stmt_2497_ack_0 : boolean;
  signal phi_stmt_2503_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5651_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5651_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5651_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5651_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5651: Block -- control-path 
    signal convTransposeC_CP_5651_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5651_elements(0) <= convTransposeC_CP_5651_start;
    convTransposeC_CP_5651_symbol <= convTransposeC_CP_5651_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2156/$entry
      -- CP-element group 0: 	 branch_block_stmt_2156/branch_block_stmt_2156__entry__
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217__entry__
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/$entry
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_update_start_
      -- 
    cr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(0), ack => type_cast_2189_inst_req_1); -- 
    cr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(0), ack => type_cast_2202_inst_req_1); -- 
    rr_5699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(0), ack => RPIPE_Block2_start_2158_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2156/merge_stmt_2489__exit__
      -- CP-element group 1: 	 branch_block_stmt_2156/assign_stmt_2515__entry__
      -- CP-element group 1: 	 branch_block_stmt_2156/assign_stmt_2515__exit__
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2156/assign_stmt_2515/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/assign_stmt_2515/$exit
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/SplitProtocol/Update/cr
      -- 
    rr_6400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(1), ack => type_cast_2288_inst_req_0); -- 
    cr_6405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(1), ack => type_cast_2288_inst_req_1); -- 
    rr_6423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(1), ack => type_cast_2295_inst_req_0); -- 
    cr_6428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(1), ack => type_cast_2295_inst_req_1); -- 
    rr_6446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(1), ack => type_cast_2302_inst_req_0); -- 
    cr_6451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(1), ack => type_cast_2302_inst_req_1); -- 
    rr_6469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(1), ack => type_cast_2308_inst_req_0); -- 
    cr_6474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(1), ack => type_cast_2308_inst_req_1); -- 
    convTransposeC_CP_5651_elements(1) <= convTransposeC_CP_5651_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_Update/cr
      -- 
    ra_5700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2158_inst_ack_0, ack => convTransposeC_CP_5651_elements(2)); -- 
    cr_5704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(2), ack => RPIPE_Block2_start_2158_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2158_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_Sample/rr
      -- 
    ca_5705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2158_inst_ack_1, ack => convTransposeC_CP_5651_elements(3)); -- 
    rr_5713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(3), ack => RPIPE_Block2_start_2161_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_Update/cr
      -- 
    ra_5714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2161_inst_ack_0, ack => convTransposeC_CP_5651_elements(4)); -- 
    cr_5718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(4), ack => RPIPE_Block2_start_2161_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2161_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_Sample/rr
      -- 
    ca_5719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2161_inst_ack_1, ack => convTransposeC_CP_5651_elements(5)); -- 
    rr_5727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(5), ack => RPIPE_Block2_start_2164_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_Update/cr
      -- 
    ra_5728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2164_inst_ack_0, ack => convTransposeC_CP_5651_elements(6)); -- 
    cr_5732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(6), ack => RPIPE_Block2_start_2164_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2164_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_Sample/rr
      -- 
    ca_5733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2164_inst_ack_1, ack => convTransposeC_CP_5651_elements(7)); -- 
    rr_5741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(7), ack => RPIPE_Block2_start_2167_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_Update/cr
      -- 
    ra_5742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2167_inst_ack_0, ack => convTransposeC_CP_5651_elements(8)); -- 
    cr_5746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(8), ack => RPIPE_Block2_start_2167_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2167_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_Sample/rr
      -- 
    ca_5747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2167_inst_ack_1, ack => convTransposeC_CP_5651_elements(9)); -- 
    rr_5755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(9), ack => RPIPE_Block2_start_2170_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_Update/cr
      -- 
    ra_5756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2170_inst_ack_0, ack => convTransposeC_CP_5651_elements(10)); -- 
    cr_5760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(10), ack => RPIPE_Block2_start_2170_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2170_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_Sample/rr
      -- 
    ca_5761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2170_inst_ack_1, ack => convTransposeC_CP_5651_elements(11)); -- 
    rr_5769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(11), ack => RPIPE_Block2_start_2173_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_Update/cr
      -- 
    ra_5770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2173_inst_ack_0, ack => convTransposeC_CP_5651_elements(12)); -- 
    cr_5774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(12), ack => RPIPE_Block2_start_2173_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2173_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_Sample/rr
      -- 
    ca_5775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2173_inst_ack_1, ack => convTransposeC_CP_5651_elements(13)); -- 
    rr_5783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(13), ack => RPIPE_Block2_start_2176_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_Update/cr
      -- 
    ra_5784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2176_inst_ack_0, ack => convTransposeC_CP_5651_elements(14)); -- 
    cr_5788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(14), ack => RPIPE_Block2_start_2176_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2176_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_Sample/rr
      -- 
    ca_5789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2176_inst_ack_1, ack => convTransposeC_CP_5651_elements(15)); -- 
    rr_5797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(15), ack => RPIPE_Block2_start_2179_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_Update/cr
      -- 
    ra_5798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2179_inst_ack_0, ack => convTransposeC_CP_5651_elements(16)); -- 
    cr_5802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(16), ack => RPIPE_Block2_start_2179_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2179_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_Sample/rr
      -- 
    ca_5803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2179_inst_ack_1, ack => convTransposeC_CP_5651_elements(17)); -- 
    rr_5811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(17), ack => RPIPE_Block2_start_2182_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_Update/cr
      -- 
    ra_5812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2182_inst_ack_0, ack => convTransposeC_CP_5651_elements(18)); -- 
    cr_5816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(18), ack => RPIPE_Block2_start_2182_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2182_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_Sample/rr
      -- 
    ca_5817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2182_inst_ack_1, ack => convTransposeC_CP_5651_elements(19)); -- 
    rr_5825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(19), ack => RPIPE_Block2_start_2185_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_Update/cr
      -- 
    ra_5826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2185_inst_ack_0, ack => convTransposeC_CP_5651_elements(20)); -- 
    cr_5830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(20), ack => RPIPE_Block2_start_2185_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2185_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_Sample/rr
      -- 
    ca_5831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2185_inst_ack_1, ack => convTransposeC_CP_5651_elements(21)); -- 
    rr_5839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(21), ack => type_cast_2189_inst_req_0); -- 
    rr_5853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(21), ack => RPIPE_Block2_start_2198_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_Sample/ra
      -- 
    ra_5840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2189_inst_ack_0, ack => convTransposeC_CP_5651_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2189_update_completed_
      -- 
    ca_5845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2189_inst_ack_1, ack => convTransposeC_CP_5651_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_update_start_
      -- 
    ra_5854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2198_inst_ack_0, ack => convTransposeC_CP_5651_elements(24)); -- 
    cr_5858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(24), ack => RPIPE_Block2_start_2198_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2198_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_Sample/rr
      -- 
    ca_5859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2198_inst_ack_1, ack => convTransposeC_CP_5651_elements(25)); -- 
    rr_5867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(25), ack => type_cast_2202_inst_req_0); -- 
    rr_5881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(25), ack => RPIPE_Block2_start_2210_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_Sample/$exit
      -- 
    ra_5868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2202_inst_ack_0, ack => convTransposeC_CP_5651_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/type_cast_2202_Update/$exit
      -- 
    ca_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2202_inst_ack_1, ack => convTransposeC_CP_5651_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_Sample/ra
      -- 
    ra_5882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2210_inst_ack_0, ack => convTransposeC_CP_5651_elements(28)); -- 
    cr_5886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(28), ack => RPIPE_Block2_start_2210_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2210_Update/$exit
      -- 
    ca_5887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2210_inst_ack_1, ack => convTransposeC_CP_5651_elements(29)); -- 
    rr_5895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(29), ack => RPIPE_Block2_start_2213_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_sample_completed_
      -- 
    ra_5896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2213_inst_ack_0, ack => convTransposeC_CP_5651_elements(30)); -- 
    cr_5900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(30), ack => RPIPE_Block2_start_2213_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2213_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_Sample/$entry
      -- 
    ca_5901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2213_inst_ack_1, ack => convTransposeC_CP_5651_elements(31)); -- 
    rr_5909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(31), ack => RPIPE_Block2_start_2216_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_update_start_
      -- 
    ra_5910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2216_inst_ack_0, ack => convTransposeC_CP_5651_elements(32)); -- 
    cr_5914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(32), ack => RPIPE_Block2_start_2216_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/RPIPE_Block2_start_2216_update_completed_
      -- 
    ca_5915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2216_inst_ack_1, ack => convTransposeC_CP_5651_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/$entry
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217__exit__
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279__entry__
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2159_to_assign_stmt_2217/$exit
      -- CP-element group 34: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_Update/cr
      -- 
    cr_5973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(34), ack => type_cast_2261_inst_req_1); -- 
    rr_5926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(34), ack => type_cast_2249_inst_req_0); -- 
    cr_5945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(34), ack => type_cast_2253_inst_req_1); -- 
    rr_5954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(34), ack => type_cast_2257_inst_req_0); -- 
    cr_5959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(34), ack => type_cast_2257_inst_req_1); -- 
    rr_5968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(34), ack => type_cast_2261_inst_req_0); -- 
    rr_5940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(34), ack => type_cast_2253_inst_req_0); -- 
    cr_5931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(34), ack => type_cast_2249_inst_req_1); -- 
    convTransposeC_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(23) & convTransposeC_CP_5651_elements(27) & convTransposeC_CP_5651_elements(33);
      gj_convTransposeC_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_sample_completed_
      -- 
    ra_5927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2249_inst_ack_0, ack => convTransposeC_CP_5651_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2249_Update/$exit
      -- 
    ca_5932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2249_inst_ack_1, ack => convTransposeC_CP_5651_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_sample_completed_
      -- 
    ra_5941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2253_inst_ack_0, ack => convTransposeC_CP_5651_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2253_update_completed_
      -- 
    ca_5946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2253_inst_ack_1, ack => convTransposeC_CP_5651_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_Sample/ra
      -- 
    ra_5955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2257_inst_ack_0, ack => convTransposeC_CP_5651_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2257_Update/ca
      -- 
    ca_5960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2257_inst_ack_1, ack => convTransposeC_CP_5651_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_sample_completed_
      -- 
    ra_5969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2261_inst_ack_0, ack => convTransposeC_CP_5651_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/type_cast_2261_update_completed_
      -- 
    ca_5974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2261_inst_ack_1, ack => convTransposeC_CP_5651_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279/$exit
      -- CP-element group 43: 	 branch_block_stmt_2156/assign_stmt_2224_to_assign_stmt_2279__exit__
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2282/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2289/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2296/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/SplitProtocol/Update/cr
      -- 
    rr_6374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(43), ack => type_cast_2306_inst_req_0); -- 
    cr_6379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(43), ack => type_cast_2306_inst_req_1); -- 
    convTransposeC_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(36) & convTransposeC_CP_5651_elements(38) & convTransposeC_CP_5651_elements(40) & convTransposeC_CP_5651_elements(42);
      gj_convTransposeC_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_Sample/$exit
      -- 
    ra_5986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2343_inst_ack_0, ack => convTransposeC_CP_5651_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_update_completed_
      -- 
    ca_5991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2343_inst_ack_1, ack => convTransposeC_CP_5651_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_sample_completed_
      -- 
    ra_6000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_0, ack => convTransposeC_CP_5651_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_Update/ca
      -- 
    ca_6005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2347_inst_ack_1, ack => convTransposeC_CP_5651_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_sample_completed_
      -- 
    ra_6014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_0, ack => convTransposeC_CP_5651_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_Update/ca
      -- 
    ca_6019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_1, ack => convTransposeC_CP_5651_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_sample_completed_
      -- 
    ra_6028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2381_inst_ack_0, ack => convTransposeC_CP_5651_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_final_index_sum_regn_Sample/req
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_index_computed_1
      -- 
    ca_6033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2381_inst_ack_1, ack => convTransposeC_CP_5651_elements(51)); -- 
    req_6058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(51), ack => array_obj_ref_2387_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_final_index_sum_regn_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_final_index_sum_regn_sample_complete
      -- 
    ack_6059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2387_index_offset_ack_0, ack => convTransposeC_CP_5651_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_request/req
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_base_plus_offset/sum_rename_ack
      -- 
    ack_6064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2387_index_offset_ack_1, ack => convTransposeC_CP_5651_elements(53)); -- 
    req_6073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(53), ack => addr_of_2388_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_request/ack
      -- CP-element group 54: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_request/$exit
      -- 
    ack_6074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2388_final_reg_ack_0, ack => convTransposeC_CP_5651_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Sample/word_access_start/word_0/rr
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_base_address_resized
      -- 
    ack_6079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2388_final_reg_ack_1, ack => convTransposeC_CP_5651_elements(55)); -- 
    rr_6112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(55), ack => ptr_deref_2392_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Sample/word_access_start/word_0/ra
      -- 
    ra_6113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2392_load_0_ack_0, ack => convTransposeC_CP_5651_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/ptr_deref_2392_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/ptr_deref_2392_Merge/merge_ack
      -- CP-element group 57: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/ptr_deref_2392_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/ptr_deref_2392_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_update_completed_
      -- 
    ca_6124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2392_load_0_ack_1, ack => convTransposeC_CP_5651_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_index_resize_1/index_resize_ack
      -- 
    req_6154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(58), ack => array_obj_ref_2410_index_offset_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(45) & convTransposeC_CP_5651_elements(47) & convTransposeC_CP_5651_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_final_index_sum_regn_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_final_index_sum_regn_sample_complete
      -- 
    ack_6155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2410_index_offset_ack_0, ack => convTransposeC_CP_5651_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_request/req
      -- 
    ack_6160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2410_index_offset_ack_1, ack => convTransposeC_CP_5651_elements(60)); -- 
    req_6169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(60), ack => addr_of_2411_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_request/ack
      -- 
    ack_6170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2411_final_reg_ack_0, ack => convTransposeC_CP_5651_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_complete/$exit
      -- 
    ack_6175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2411_final_reg_ack_1, ack => convTransposeC_CP_5651_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/ptr_deref_2414_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/ptr_deref_2414_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/ptr_deref_2414_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/ptr_deref_2414_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/word_access_start/word_0/rr
      -- 
    rr_6213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(63), ack => ptr_deref_2414_store_0_req_0); -- 
    convTransposeC_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(57) & convTransposeC_CP_5651_elements(62);
      gj_convTransposeC_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Sample/word_access_start/word_0/ra
      -- 
    ra_6214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2414_store_0_ack_0, ack => convTransposeC_CP_5651_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Update/word_access_complete/word_0/ca
      -- 
    ca_6225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2414_store_0_ack_1, ack => convTransposeC_CP_5651_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_Sample/ra
      -- 
    ra_6234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2419_inst_ack_0, ack => convTransposeC_CP_5651_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_Update/ca
      -- 
    ca_6239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2419_inst_ack_1, ack => convTransposeC_CP_5651_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/$exit
      -- CP-element group 68: 	 branch_block_stmt_2156/R_cmp_2433_place
      -- CP-element group 68: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431__exit__
      -- CP-element group 68: 	 branch_block_stmt_2156/if_stmt_2432__entry__
      -- CP-element group 68: 	 branch_block_stmt_2156/if_stmt_2432_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2156/if_stmt_2432_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_2156/if_stmt_2432_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_2156/if_stmt_2432_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_2156/if_stmt_2432_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2156/if_stmt_2432_else_link/$entry
      -- 
    branch_req_6247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(68), ack => if_stmt_2432_branch_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(52) & convTransposeC_CP_5651_elements(59) & convTransposeC_CP_5651_elements(65) & convTransposeC_CP_5651_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_2156/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_2156/merge_stmt_2438__exit__
      -- CP-element group 69: 	 branch_block_stmt_2156/assign_stmt_2444__entry__
      -- CP-element group 69: 	 branch_block_stmt_2156/assign_stmt_2444__exit__
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133
      -- CP-element group 69: 	 branch_block_stmt_2156/if_stmt_2432_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_2156/if_stmt_2432_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_2156/assign_stmt_2444/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/assign_stmt_2444/$exit
      -- CP-element group 69: 	 branch_block_stmt_2156/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_2156/merge_stmt_2438_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_2156/merge_stmt_2438_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/merge_stmt_2438_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_2156/merge_stmt_2438_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2432_branch_ack_1, ack => convTransposeC_CP_5651_elements(69)); -- 
    rr_6584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(69), ack => type_cast_2493_inst_req_0); -- 
    cr_6589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(69), ack => type_cast_2493_inst_req_1); -- 
    rr_6607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(69), ack => type_cast_2502_inst_req_0); -- 
    cr_6612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(69), ack => type_cast_2502_inst_req_1); -- 
    rr_6630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(69), ack => type_cast_2508_inst_req_0); -- 
    cr_6635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(69), ack => type_cast_2508_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_2156/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_2156/merge_stmt_2446__exit__
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482__entry__
      -- CP-element group 70: 	 branch_block_stmt_2156/if_stmt_2432_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_2156/if_stmt_2432_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/$entry
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2156/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2156/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2156/merge_stmt_2446_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2156/merge_stmt_2446_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2156/merge_stmt_2446_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2156/merge_stmt_2446_PhiAck/dummy
      -- 
    else_choice_transition_6256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2432_branch_ack_0, ack => convTransposeC_CP_5651_elements(70)); -- 
    rr_6272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(70), ack => type_cast_2460_inst_req_0); -- 
    cr_6277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(70), ack => type_cast_2460_inst_req_1); -- 
    cr_6291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(70), ack => type_cast_2476_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_Sample/ra
      -- 
    ra_6273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_0, ack => convTransposeC_CP_5651_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2460_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_Sample/rr
      -- 
    ca_6278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_1, ack => convTransposeC_CP_5651_elements(72)); -- 
    rr_6286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(72), ack => type_cast_2476_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_Sample/ra
      -- 
    ra_6287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2476_inst_ack_0, ack => convTransposeC_CP_5651_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_2156/R_cmp122_2484_place
      -- CP-element group 74: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482__exit__
      -- CP-element group 74: 	 branch_block_stmt_2156/if_stmt_2483__entry__
      -- CP-element group 74: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/$exit
      -- CP-element group 74: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2156/assign_stmt_2452_to_assign_stmt_2482/type_cast_2476_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_2156/if_stmt_2483_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2156/if_stmt_2483_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_2156/if_stmt_2483_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_2156/if_stmt_2483_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_2156/if_stmt_2483_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2156/if_stmt_2483_else_link/$entry
      -- 
    ca_6292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2476_inst_ack_1, ack => convTransposeC_CP_5651_elements(74)); -- 
    branch_req_6300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(74), ack => if_stmt_2483_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_2156/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_2156/merge_stmt_2517__exit__
      -- CP-element group 75: 	 branch_block_stmt_2156/assign_stmt_2522__entry__
      -- CP-element group 75: 	 branch_block_stmt_2156/if_stmt_2483_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_2156/if_stmt_2483_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_2156/assign_stmt_2522/$entry
      -- CP-element group 75: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_2156/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2156/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_2156/merge_stmt_2517_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_2156/merge_stmt_2517_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_2156/merge_stmt_2517_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2156/merge_stmt_2517_PhiAck/dummy
      -- 
    if_choice_transition_6305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2483_branch_ack_1, ack => convTransposeC_CP_5651_elements(75)); -- 
    req_6325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(75), ack => WPIPE_Block2_done_2519_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133
      -- CP-element group 76: 	 branch_block_stmt_2156/if_stmt_2483_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_2156/if_stmt_2483_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2490/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2483_branch_ack_0, ack => convTransposeC_CP_5651_elements(76)); -- 
    rr_6535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(76), ack => type_cast_2500_inst_req_0); -- 
    cr_6540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(76), ack => type_cast_2500_inst_req_1); -- 
    rr_6558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(76), ack => type_cast_2506_inst_req_0); -- 
    cr_6563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(76), ack => type_cast_2506_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_Update/req
      -- 
    ack_6326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2519_inst_ack_0, ack => convTransposeC_CP_5651_elements(77)); -- 
    req_6330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(77), ack => WPIPE_Block2_done_2519_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_2156/$exit
      -- CP-element group 78: 	 branch_block_stmt_2156/branch_block_stmt_2156__exit__
      -- CP-element group 78: 	 branch_block_stmt_2156/assign_stmt_2522__exit__
      -- CP-element group 78: 	 branch_block_stmt_2156/return__
      -- CP-element group 78: 	 branch_block_stmt_2156/merge_stmt_2524__exit__
      -- CP-element group 78: 	 branch_block_stmt_2156/assign_stmt_2522/$exit
      -- CP-element group 78: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2156/assign_stmt_2522/WPIPE_Block2_done_2519_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_2156/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2156/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2156/merge_stmt_2524_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2156/merge_stmt_2524_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2156/merge_stmt_2524_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2156/merge_stmt_2524_PhiAck/dummy
      -- 
    ack_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2519_inst_ack_1, ack => convTransposeC_CP_5651_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	85 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2282/$exit
      -- CP-element group 79: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2286_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_req
      -- 
    phi_stmt_2282_req_6342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2282_req_6342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(79), ack => phi_stmt_2282_req_0); -- 
    -- Element group convTransposeC_CP_5651_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeC_CP_5651_elements(43), ack => convTransposeC_CP_5651_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	85 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2289/$exit
      -- CP-element group 80: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2293_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_req
      -- 
    phi_stmt_2289_req_6350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2289_req_6350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(80), ack => phi_stmt_2289_req_0); -- 
    -- Element group convTransposeC_CP_5651_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeC_CP_5651_elements(43), ack => convTransposeC_CP_5651_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2296/$exit
      -- CP-element group 81: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2300_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_req
      -- 
    phi_stmt_2296_req_6358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2296_req_6358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(81), ack => phi_stmt_2296_req_0); -- 
    -- Element group convTransposeC_CP_5651_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeC_CP_5651_elements(43), ack => convTransposeC_CP_5651_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/SplitProtocol/Sample/ra
      -- 
    ra_6375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2306_inst_ack_0, ack => convTransposeC_CP_5651_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/SplitProtocol/Update/ca
      -- 
    ca_6380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2306_inst_ack_1, ack => convTransposeC_CP_5651_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/$exit
      -- CP-element group 84: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/$exit
      -- CP-element group 84: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2306/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_req
      -- 
    phi_stmt_2303_req_6381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2303_req_6381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(84), ack => phi_stmt_2303_req_0); -- 
    convTransposeC_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(82) & convTransposeC_CP_5651_elements(83);
      gj_convTransposeC_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: 	80 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2156/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(79) & convTransposeC_CP_5651_elements(80) & convTransposeC_CP_5651_elements(81) & convTransposeC_CP_5651_elements(84);
      gj_convTransposeC_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Sample/ra
      -- 
    ra_6401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2288_inst_ack_0, ack => convTransposeC_CP_5651_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/Update/ca
      -- 
    ca_6406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2288_inst_ack_1, ack => convTransposeC_CP_5651_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/$exit
      -- CP-element group 88: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/$exit
      -- CP-element group 88: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_sources/type_cast_2288/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2282/phi_stmt_2282_req
      -- 
    phi_stmt_2282_req_6407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2282_req_6407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(88), ack => phi_stmt_2282_req_1); -- 
    convTransposeC_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(86) & convTransposeC_CP_5651_elements(87);
      gj_convTransposeC_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Sample/ra
      -- 
    ra_6424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2295_inst_ack_0, ack => convTransposeC_CP_5651_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/Update/ca
      -- 
    ca_6429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2295_inst_ack_1, ack => convTransposeC_CP_5651_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/$exit
      -- CP-element group 91: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/$exit
      -- CP-element group 91: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_sources/type_cast_2295/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2289/phi_stmt_2289_req
      -- 
    phi_stmt_2289_req_6430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2289_req_6430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(91), ack => phi_stmt_2289_req_1); -- 
    convTransposeC_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(89) & convTransposeC_CP_5651_elements(90);
      gj_convTransposeC_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/SplitProtocol/Sample/ra
      -- 
    ra_6447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2302_inst_ack_0, ack => convTransposeC_CP_5651_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/SplitProtocol/Update/ca
      -- 
    ca_6452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2302_inst_ack_1, ack => convTransposeC_CP_5651_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/$exit
      -- CP-element group 94: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/$exit
      -- CP-element group 94: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_sources/type_cast_2302/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2296/phi_stmt_2296_req
      -- 
    phi_stmt_2296_req_6453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2296_req_6453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(94), ack => phi_stmt_2296_req_1); -- 
    convTransposeC_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(92) & convTransposeC_CP_5651_elements(93);
      gj_convTransposeC_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/SplitProtocol/Sample/ra
      -- 
    ra_6470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2308_inst_ack_0, ack => convTransposeC_CP_5651_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/SplitProtocol/Update/ca
      -- 
    ca_6475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2308_inst_ack_1, ack => convTransposeC_CP_5651_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/$exit
      -- CP-element group 97: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/$exit
      -- CP-element group 97: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_sources/type_cast_2308/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2303/phi_stmt_2303_req
      -- 
    phi_stmt_2303_req_6476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2303_req_6476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(97), ack => phi_stmt_2303_req_1); -- 
    convTransposeC_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(95) & convTransposeC_CP_5651_elements(96);
      gj_convTransposeC_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2156/ifx_xend133_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(88) & convTransposeC_CP_5651_elements(91) & convTransposeC_CP_5651_elements(94) & convTransposeC_CP_5651_elements(97);
      gj_convTransposeC_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2156/merge_stmt_2281_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_2156/merge_stmt_2281_PhiAck/$entry
      -- 
    convTransposeC_CP_5651_elements(99) <= OrReduce(convTransposeC_CP_5651_elements(85) & convTransposeC_CP_5651_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2156/merge_stmt_2281_PhiAck/phi_stmt_2282_ack
      -- 
    phi_stmt_2282_ack_6481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2282_ack_0, ack => convTransposeC_CP_5651_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2156/merge_stmt_2281_PhiAck/phi_stmt_2289_ack
      -- 
    phi_stmt_2289_ack_6482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2289_ack_0, ack => convTransposeC_CP_5651_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2156/merge_stmt_2281_PhiAck/phi_stmt_2296_ack
      -- 
    phi_stmt_2296_ack_6483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2296_ack_0, ack => convTransposeC_CP_5651_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2156/merge_stmt_2281_PhiAck/phi_stmt_2303_ack
      -- 
    phi_stmt_2303_ack_6484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2303_ack_0, ack => convTransposeC_CP_5651_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2387_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2347_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2392_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/array_obj_ref_2410_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2381_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2343_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2388_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/addr_of_2411_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2351_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2156/merge_stmt_2281__exit__
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431__entry__
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/ptr_deref_2414_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2156/assign_stmt_2315_to_assign_stmt_2431/type_cast_2419_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2156/merge_stmt_2281_PhiAck/$exit
      -- 
    cr_5990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => type_cast_2343_inst_req_1); -- 
    cr_6004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => type_cast_2347_inst_req_1); -- 
    rr_5999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => type_cast_2347_inst_req_0); -- 
    rr_6013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => type_cast_2351_inst_req_0); -- 
    rr_6027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => type_cast_2381_inst_req_0); -- 
    cr_6032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => type_cast_2381_inst_req_1); -- 
    req_6063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => array_obj_ref_2387_index_offset_req_1); -- 
    rr_5985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => type_cast_2343_inst_req_0); -- 
    req_6159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => array_obj_ref_2410_index_offset_req_1); -- 
    cr_6123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => ptr_deref_2392_load_0_req_1); -- 
    req_6078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => addr_of_2388_final_reg_req_1); -- 
    req_6174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => addr_of_2411_final_reg_req_1); -- 
    cr_6018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => type_cast_2351_inst_req_1); -- 
    cr_6224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => ptr_deref_2414_store_0_req_1); -- 
    rr_6233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => type_cast_2419_inst_req_0); -- 
    cr_6238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(104), ack => type_cast_2419_inst_req_1); -- 
    convTransposeC_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(100) & convTransposeC_CP_5651_elements(101) & convTransposeC_CP_5651_elements(102) & convTransposeC_CP_5651_elements(103);
      gj_convTransposeC_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  output  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2490/$exit
      -- CP-element group 105: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2496_konst_delay_trans
      -- CP-element group 105: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_req
      -- 
    phi_stmt_2490_req_6519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2490_req_6519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(105), ack => phi_stmt_2490_req_1); -- 
    -- Element group convTransposeC_CP_5651_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => convTransposeC_CP_5651_elements(76), ack => convTransposeC_CP_5651_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/SplitProtocol/Sample/ra
      -- 
    ra_6536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2500_inst_ack_0, ack => convTransposeC_CP_5651_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/SplitProtocol/Update/ca
      -- 
    ca_6541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2500_inst_ack_1, ack => convTransposeC_CP_5651_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/$exit
      -- CP-element group 108: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/$exit
      -- CP-element group 108: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2500/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_req
      -- 
    phi_stmt_2497_req_6542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2497_req_6542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(108), ack => phi_stmt_2497_req_0); -- 
    convTransposeC_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(106) & convTransposeC_CP_5651_elements(107);
      gj_convTransposeC_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Sample/ra
      -- 
    ra_6559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2506_inst_ack_0, ack => convTransposeC_CP_5651_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/Update/ca
      -- 
    ca_6564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2506_inst_ack_1, ack => convTransposeC_CP_5651_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/$exit
      -- CP-element group 111: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/$exit
      -- CP-element group 111: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2506/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_req
      -- 
    phi_stmt_2503_req_6565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2503_req_6565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(111), ack => phi_stmt_2503_req_0); -- 
    convTransposeC_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(109) & convTransposeC_CP_5651_elements(110);
      gj_convTransposeC_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2156/ifx_xelse_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(105) & convTransposeC_CP_5651_elements(108) & convTransposeC_CP_5651_elements(111);
      gj_convTransposeC_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/SplitProtocol/Sample/ra
      -- 
    ra_6585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2493_inst_ack_0, ack => convTransposeC_CP_5651_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/SplitProtocol/Update/ca
      -- 
    ca_6590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2493_inst_ack_1, ack => convTransposeC_CP_5651_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/$exit
      -- CP-element group 115: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/$exit
      -- CP-element group 115: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_sources/type_cast_2493/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2490/phi_stmt_2490_req
      -- 
    phi_stmt_2490_req_6591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2490_req_6591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(115), ack => phi_stmt_2490_req_0); -- 
    convTransposeC_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(113) & convTransposeC_CP_5651_elements(114);
      gj_convTransposeC_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/SplitProtocol/Sample/ra
      -- 
    ra_6608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2502_inst_ack_0, ack => convTransposeC_CP_5651_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/SplitProtocol/Update/ca
      -- 
    ca_6613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2502_inst_ack_1, ack => convTransposeC_CP_5651_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/$exit
      -- CP-element group 118: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/$exit
      -- CP-element group 118: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_sources/type_cast_2502/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2497/phi_stmt_2497_req
      -- 
    phi_stmt_2497_req_6614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2497_req_6614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(118), ack => phi_stmt_2497_req_1); -- 
    convTransposeC_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(116) & convTransposeC_CP_5651_elements(117);
      gj_convTransposeC_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Sample/ra
      -- 
    ra_6631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_0, ack => convTransposeC_CP_5651_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/Update/ca
      -- 
    ca_6636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_1, ack => convTransposeC_CP_5651_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/$exit
      -- CP-element group 121: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/$exit
      -- CP-element group 121: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_sources/type_cast_2508/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2503/phi_stmt_2503_req
      -- 
    phi_stmt_2503_req_6637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2503_req_6637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5651_elements(121), ack => phi_stmt_2503_req_1); -- 
    convTransposeC_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(119) & convTransposeC_CP_5651_elements(120);
      gj_convTransposeC_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2156/ifx_xthen_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(115) & convTransposeC_CP_5651_elements(118) & convTransposeC_CP_5651_elements(121);
      gj_convTransposeC_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2156/merge_stmt_2489_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_2156/merge_stmt_2489_PhiAck/$entry
      -- 
    convTransposeC_CP_5651_elements(123) <= OrReduce(convTransposeC_CP_5651_elements(112) & convTransposeC_CP_5651_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2156/merge_stmt_2489_PhiAck/phi_stmt_2490_ack
      -- 
    phi_stmt_2490_ack_6642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2490_ack_0, ack => convTransposeC_CP_5651_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2156/merge_stmt_2489_PhiAck/phi_stmt_2497_ack
      -- 
    phi_stmt_2497_ack_6643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2497_ack_0, ack => convTransposeC_CP_5651_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2156/merge_stmt_2489_PhiAck/phi_stmt_2503_ack
      -- 
    phi_stmt_2503_ack_6644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2503_ack_0, ack => convTransposeC_CP_5651_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2156/merge_stmt_2489_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5651_elements(124) & convTransposeC_CP_5651_elements(125) & convTransposeC_CP_5651_elements(126);
      gj_convTransposeC_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5651_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2409_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2409_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2386_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2386_scaled : std_logic_vector(13 downto 0);
    signal add121_2279 : std_logic_vector(31 downto 0);
    signal add45_2230 : std_logic_vector(15 downto 0);
    signal add58_2241 : std_logic_vector(15 downto 0);
    signal add77_2362 : std_logic_vector(63 downto 0);
    signal add79_2372 : std_logic_vector(63 downto 0);
    signal add91_2426 : std_logic_vector(31 downto 0);
    signal add98_2444 : std_logic_vector(15 downto 0);
    signal add_2208 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2320 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2387_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2387_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2387_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2387_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2387_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2387_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2410_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2410_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2410_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2410_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2410_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2410_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2389 : std_logic_vector(31 downto 0);
    signal arrayidx87_2412 : std_logic_vector(31 downto 0);
    signal call11_2177 : std_logic_vector(15 downto 0);
    signal call13_2180 : std_logic_vector(15 downto 0);
    signal call14_2183 : std_logic_vector(15 downto 0);
    signal call15_2186 : std_logic_vector(15 downto 0);
    signal call16_2199 : std_logic_vector(15 downto 0);
    signal call18_2211 : std_logic_vector(15 downto 0);
    signal call1_2162 : std_logic_vector(15 downto 0);
    signal call20_2214 : std_logic_vector(15 downto 0);
    signal call22_2217 : std_logic_vector(15 downto 0);
    signal call3_2165 : std_logic_vector(15 downto 0);
    signal call5_2168 : std_logic_vector(15 downto 0);
    signal call7_2171 : std_logic_vector(15 downto 0);
    signal call9_2174 : std_logic_vector(15 downto 0);
    signal call_2159 : std_logic_vector(15 downto 0);
    signal cmp106_2457 : std_logic_vector(0 downto 0);
    signal cmp122_2482 : std_logic_vector(0 downto 0);
    signal cmp_2431 : std_logic_vector(0 downto 0);
    signal conv112_2477 : std_logic_vector(31 downto 0);
    signal conv115_2262 : std_logic_vector(31 downto 0);
    signal conv17_2203 : std_logic_vector(31 downto 0);
    signal conv65_2344 : std_logic_vector(63 downto 0);
    signal conv68_2250 : std_logic_vector(63 downto 0);
    signal conv70_2348 : std_logic_vector(63 downto 0);
    signal conv73_2254 : std_logic_vector(63 downto 0);
    signal conv75_2352 : std_logic_vector(63 downto 0);
    signal conv90_2420 : std_logic_vector(31 downto 0);
    signal conv94_2258 : std_logic_vector(31 downto 0);
    signal conv_2190 : std_logic_vector(31 downto 0);
    signal idxprom86_2405 : std_logic_vector(63 downto 0);
    signal idxprom_2382 : std_logic_vector(63 downto 0);
    signal inc110_2461 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2466 : std_logic_vector(15 downto 0);
    signal inc_2452 : std_logic_vector(15 downto 0);
    signal indvar_2282 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2515 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2503 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2303 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2497 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2296 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2473 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2490 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2289 : std_logic_vector(15 downto 0);
    signal mul54_2335 : std_logic_vector(15 downto 0);
    signal mul76_2357 : std_logic_vector(63 downto 0);
    signal mul78_2367 : std_logic_vector(63 downto 0);
    signal mul_2325 : std_logic_vector(15 downto 0);
    signal ptr_deref_2392_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2392_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2392_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2392_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2392_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2414_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2414_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2414_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2414_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2414_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2414_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2196 : std_logic_vector(31 downto 0);
    signal shr116137_2268 : std_logic_vector(31 downto 0);
    signal shr120138_2274 : std_logic_vector(31 downto 0);
    signal shr136_2224 : std_logic_vector(15 downto 0);
    signal shr81_2378 : std_logic_vector(31 downto 0);
    signal shr85_2399 : std_logic_vector(63 downto 0);
    signal sub48_2330 : std_logic_vector(15 downto 0);
    signal sub61_2246 : std_logic_vector(15 downto 0);
    signal sub62_2340 : std_logic_vector(15 downto 0);
    signal sub_2235 : std_logic_vector(15 downto 0);
    signal tmp1_2315 : std_logic_vector(31 downto 0);
    signal tmp83_2393 : std_logic_vector(63 downto 0);
    signal type_cast_2194_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2222_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2228_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2239_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2266_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2272_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2286_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2288_wire : std_logic_vector(31 downto 0);
    signal type_cast_2293_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2295_wire : std_logic_vector(15 downto 0);
    signal type_cast_2300_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2302_wire : std_logic_vector(15 downto 0);
    signal type_cast_2306_wire : std_logic_vector(15 downto 0);
    signal type_cast_2308_wire : std_logic_vector(15 downto 0);
    signal type_cast_2313_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2376_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2397_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2403_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2424_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2442_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2450_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2470_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2493_wire : std_logic_vector(15 downto 0);
    signal type_cast_2496_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2500_wire : std_logic_vector(15 downto 0);
    signal type_cast_2502_wire : std_logic_vector(15 downto 0);
    signal type_cast_2506_wire : std_logic_vector(15 downto 0);
    signal type_cast_2508_wire : std_logic_vector(15 downto 0);
    signal type_cast_2513_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2521_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2387_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2387_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2387_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2387_resized_base_address <= "00000000000000";
    array_obj_ref_2410_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2410_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2410_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2410_resized_base_address <= "00000000000000";
    ptr_deref_2392_word_offset_0 <= "00000000000000";
    ptr_deref_2414_word_offset_0 <= "00000000000000";
    type_cast_2194_wire_constant <= "00000000000000000000000000010000";
    type_cast_2222_wire_constant <= "0000000000000001";
    type_cast_2228_wire_constant <= "1111111111111111";
    type_cast_2239_wire_constant <= "1111111111111111";
    type_cast_2266_wire_constant <= "00000000000000000000000000000010";
    type_cast_2272_wire_constant <= "00000000000000000000000000000001";
    type_cast_2286_wire_constant <= "00000000000000000000000000000000";
    type_cast_2293_wire_constant <= "0000000000000000";
    type_cast_2300_wire_constant <= "0000000000000000";
    type_cast_2313_wire_constant <= "00000000000000000000000000000100";
    type_cast_2376_wire_constant <= "00000000000000000000000000000010";
    type_cast_2397_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2403_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2424_wire_constant <= "00000000000000000000000000000100";
    type_cast_2442_wire_constant <= "0000000000000100";
    type_cast_2450_wire_constant <= "0000000000000001";
    type_cast_2470_wire_constant <= "0000000000000000";
    type_cast_2496_wire_constant <= "0000000000000000";
    type_cast_2513_wire_constant <= "00000000000000000000000000000001";
    type_cast_2521_wire_constant <= "0000000000000001";
    phi_stmt_2282: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2286_wire_constant & type_cast_2288_wire;
      req <= phi_stmt_2282_req_0 & phi_stmt_2282_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2282",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2282_ack_0,
          idata => idata,
          odata => indvar_2282,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2282
    phi_stmt_2289: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2293_wire_constant & type_cast_2295_wire;
      req <= phi_stmt_2289_req_0 & phi_stmt_2289_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2289",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2289_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2289,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2289
    phi_stmt_2296: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2300_wire_constant & type_cast_2302_wire;
      req <= phi_stmt_2296_req_0 & phi_stmt_2296_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2296",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2296_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2296,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2296
    phi_stmt_2303: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2306_wire & type_cast_2308_wire;
      req <= phi_stmt_2303_req_0 & phi_stmt_2303_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2303",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2303_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2303,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2303
    phi_stmt_2490: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2493_wire & type_cast_2496_wire_constant;
      req <= phi_stmt_2490_req_0 & phi_stmt_2490_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2490",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2490_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2490,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2490
    phi_stmt_2497: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2500_wire & type_cast_2502_wire;
      req <= phi_stmt_2497_req_0 & phi_stmt_2497_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2497",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2497_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2497,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2497
    phi_stmt_2503: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2506_wire & type_cast_2508_wire;
      req <= phi_stmt_2503_req_0 & phi_stmt_2503_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2503",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2503_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2503,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2503
    -- flow-through select operator MUX_2472_inst
    input_dim1x_x2_2473 <= type_cast_2470_wire_constant when (cmp106_2457(0) /=  '0') else inc_2452;
    addr_of_2388_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2388_final_reg_req_0;
      addr_of_2388_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2388_final_reg_req_1;
      addr_of_2388_final_reg_ack_1<= rack(0);
      addr_of_2388_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2388_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2387_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2411_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2411_final_reg_req_0;
      addr_of_2411_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2411_final_reg_req_1;
      addr_of_2411_final_reg_ack_1<= rack(0);
      addr_of_2411_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2411_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2410_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2412,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2189_inst_req_0;
      type_cast_2189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2189_inst_req_1;
      type_cast_2189_inst_ack_1<= rack(0);
      type_cast_2189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2190,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2202_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2202_inst_req_0;
      type_cast_2202_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2202_inst_req_1;
      type_cast_2202_inst_ack_1<= rack(0);
      type_cast_2202_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2202_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2203,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2249_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2249_inst_req_0;
      type_cast_2249_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2249_inst_req_1;
      type_cast_2249_inst_ack_1<= rack(0);
      type_cast_2249_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2249_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2250,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2253_inst_req_0;
      type_cast_2253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2253_inst_req_1;
      type_cast_2253_inst_ack_1<= rack(0);
      type_cast_2253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2214,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2257_inst_req_0;
      type_cast_2257_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2257_inst_req_1;
      type_cast_2257_inst_ack_1<= rack(0);
      type_cast_2257_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2257_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2258,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2261_inst_req_0;
      type_cast_2261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2261_inst_req_1;
      type_cast_2261_inst_ack_1<= rack(0);
      type_cast_2261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2159,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_2262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2288_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2288_inst_req_0;
      type_cast_2288_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2288_inst_req_1;
      type_cast_2288_inst_ack_1<= rack(0);
      type_cast_2288_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2288_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2288_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2295_inst_req_0;
      type_cast_2295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2295_inst_req_1;
      type_cast_2295_inst_ack_1<= rack(0);
      type_cast_2295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2490,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2295_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2302_inst_req_0;
      type_cast_2302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2302_inst_req_1;
      type_cast_2302_inst_ack_1<= rack(0);
      type_cast_2302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2497,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2302_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2306_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2306_inst_req_0;
      type_cast_2306_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2306_inst_req_1;
      type_cast_2306_inst_ack_1<= rack(0);
      type_cast_2306_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2306_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr136_2224,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2306_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2308_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2308_inst_req_0;
      type_cast_2308_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2308_inst_req_1;
      type_cast_2308_inst_ack_1<= rack(0);
      type_cast_2308_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2308_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2503,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2308_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2343_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2343_inst_req_0;
      type_cast_2343_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2343_inst_req_1;
      type_cast_2343_inst_ack_1<= rack(0);
      type_cast_2343_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2343_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2344,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2347_inst_req_0;
      type_cast_2347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2347_inst_req_1;
      type_cast_2347_inst_ack_1<= rack(0);
      type_cast_2347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2340,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2348,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2351_inst_req_0;
      type_cast_2351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2351_inst_req_1;
      type_cast_2351_inst_ack_1<= rack(0);
      type_cast_2351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2330,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2381_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2381_inst_req_0;
      type_cast_2381_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2381_inst_req_1;
      type_cast_2381_inst_ack_1<= rack(0);
      type_cast_2381_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2381_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2382,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2419_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2419_inst_req_0;
      type_cast_2419_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2419_inst_req_1;
      type_cast_2419_inst_ack_1<= rack(0);
      type_cast_2419_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2419_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2420,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2460_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2460_inst_req_0;
      type_cast_2460_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2460_inst_req_1;
      type_cast_2460_inst_ack_1<= rack(0);
      type_cast_2460_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2460_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2457,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2461,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2476_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2476_inst_req_0;
      type_cast_2476_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2476_inst_req_1;
      type_cast_2476_inst_ack_1<= rack(0);
      type_cast_2476_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2476_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2466,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2477,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2493_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2493_inst_req_0;
      type_cast_2493_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2493_inst_req_1;
      type_cast_2493_inst_ack_1<= rack(0);
      type_cast_2493_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2493_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2444,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2493_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2500_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2500_inst_req_0;
      type_cast_2500_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2500_inst_req_1;
      type_cast_2500_inst_ack_1<= rack(0);
      type_cast_2500_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2500_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2473,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2500_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2502_inst_req_0;
      type_cast_2502_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2502_inst_req_1;
      type_cast_2502_inst_ack_1<= rack(0);
      type_cast_2502_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2502_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2296,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2502_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2506_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2506_inst_req_0;
      type_cast_2506_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2506_inst_req_1;
      type_cast_2506_inst_ack_1<= rack(0);
      type_cast_2506_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2506_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2466,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2506_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2508_inst_req_0;
      type_cast_2508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2508_inst_req_1;
      type_cast_2508_inst_ack_1<= rack(0);
      type_cast_2508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2303,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2508_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2387_index_1_rename
    process(R_idxprom_2386_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2386_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2386_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2387_index_1_resize
    process(idxprom_2382) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2382;
      ov := iv(13 downto 0);
      R_idxprom_2386_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2387_root_address_inst
    process(array_obj_ref_2387_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2387_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2387_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2410_index_1_rename
    process(R_idxprom86_2409_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2409_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2409_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2410_index_1_resize
    process(idxprom86_2405) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2405;
      ov := iv(13 downto 0);
      R_idxprom86_2409_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2410_root_address_inst
    process(array_obj_ref_2410_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2410_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2410_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2392_addr_0
    process(ptr_deref_2392_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2392_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2392_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2392_base_resize
    process(arrayidx82_2389) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2389;
      ov := iv(13 downto 0);
      ptr_deref_2392_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2392_gather_scatter
    process(ptr_deref_2392_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2392_data_0;
      ov(63 downto 0) := iv;
      tmp83_2393 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2392_root_address_inst
    process(ptr_deref_2392_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2392_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2392_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2414_addr_0
    process(ptr_deref_2414_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2414_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2414_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2414_base_resize
    process(arrayidx87_2412) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2412;
      ov := iv(13 downto 0);
      ptr_deref_2414_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2414_gather_scatter
    process(tmp83_2393) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2393;
      ov(63 downto 0) := iv;
      ptr_deref_2414_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2414_root_address_inst
    process(ptr_deref_2414_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2414_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2414_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2432_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2431;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2432_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2432_branch_req_0,
          ack0 => if_stmt_2432_branch_ack_0,
          ack1 => if_stmt_2432_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2483_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp122_2482;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2483_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2483_branch_req_0,
          ack0 => if_stmt_2483_branch_ack_0,
          ack1 => if_stmt_2483_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2229_inst
    process(call7_2171) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2171, type_cast_2228_wire_constant, tmp_var);
      add45_2230 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2240_inst
    process(call9_2174) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2174, type_cast_2239_wire_constant, tmp_var);
      add58_2241 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2329_inst
    process(sub_2235, mul_2325) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2235, mul_2325, tmp_var);
      sub48_2330 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2339_inst
    process(sub61_2246, mul54_2335) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_2246, mul54_2335, tmp_var);
      sub62_2340 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2443_inst
    process(input_dim2x_x1_2289) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2289, type_cast_2442_wire_constant, tmp_var);
      add98_2444 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2451_inst
    process(input_dim1x_x1_2296) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2296, type_cast_2450_wire_constant, tmp_var);
      inc_2452 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2465_inst
    process(inc110_2461, input_dim0x_x2_2303) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2461, input_dim0x_x2_2303, tmp_var);
      inc110x_xinput_dim0x_x2_2466 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2278_inst
    process(shr116137_2268, shr120138_2274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr116137_2268, shr120138_2274, tmp_var);
      add121_2279 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2319_inst
    process(add_2208, tmp1_2315) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2208, tmp1_2315, tmp_var);
      add_src_0x_x0_2320 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2425_inst
    process(conv90_2420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2420, type_cast_2424_wire_constant, tmp_var);
      add91_2426 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2514_inst
    process(indvar_2282) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2282, type_cast_2513_wire_constant, tmp_var);
      indvarx_xnext_2515 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2361_inst
    process(mul76_2357, conv70_2348) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2357, conv70_2348, tmp_var);
      add77_2362 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2371_inst
    process(mul78_2367, conv65_2344) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2367, conv65_2344, tmp_var);
      add79_2372 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2404_inst
    process(shr85_2399) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2399, type_cast_2403_wire_constant, tmp_var);
      idxprom86_2405 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2456_inst
    process(inc_2452, call1_2162) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2452, call1_2162, tmp_var);
      cmp106_2457 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2481_inst
    process(conv112_2477, add121_2279) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2477, add121_2279, tmp_var);
      cmp122_2482 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2223_inst
    process(call_2159) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2159, type_cast_2222_wire_constant, tmp_var);
      shr136_2224 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2267_inst
    process(conv115_2262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2262, type_cast_2266_wire_constant, tmp_var);
      shr116137_2268 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2273_inst
    process(conv115_2262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2262, type_cast_2272_wire_constant, tmp_var);
      shr120138_2274 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2377_inst
    process(add_src_0x_x0_2320) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2320, type_cast_2376_wire_constant, tmp_var);
      shr81_2378 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2398_inst
    process(add79_2372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2372, type_cast_2397_wire_constant, tmp_var);
      shr85_2399 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2324_inst
    process(input_dim0x_x2_2303, call13_2180) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2303, call13_2180, tmp_var);
      mul_2325 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2334_inst
    process(input_dim1x_x1_2296, call13_2180) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2296, call13_2180, tmp_var);
      mul54_2335 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2314_inst
    process(indvar_2282) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2282, type_cast_2313_wire_constant, tmp_var);
      tmp1_2315 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2356_inst
    process(conv75_2352, conv73_2254) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2352, conv73_2254, tmp_var);
      mul76_2357 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2366_inst
    process(add77_2362, conv68_2250) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2362, conv68_2250, tmp_var);
      mul78_2367 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2207_inst
    process(shl_2196, conv17_2203) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2196, conv17_2203, tmp_var);
      add_2208 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2195_inst
    process(conv_2190) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2190, type_cast_2194_wire_constant, tmp_var);
      shl_2196 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2234_inst
    process(add45_2230, call14_2183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_2230, call14_2183, tmp_var);
      sub_2235 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2245_inst
    process(add58_2241, call14_2183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_2241, call14_2183, tmp_var);
      sub61_2246 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2430_inst
    process(add91_2426, conv94_2258) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2426, conv94_2258, tmp_var);
      cmp_2431 <= tmp_var; --
    end process;
    -- shared split operator group (31) : array_obj_ref_2387_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2386_scaled;
      array_obj_ref_2387_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2387_index_offset_req_0;
      array_obj_ref_2387_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2387_index_offset_req_1;
      array_obj_ref_2387_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_2410_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2409_scaled;
      array_obj_ref_2410_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2410_index_offset_req_0;
      array_obj_ref_2410_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2410_index_offset_req_1;
      array_obj_ref_2410_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared load operator group (0) : ptr_deref_2392_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2392_load_0_req_0;
      ptr_deref_2392_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2392_load_0_req_1;
      ptr_deref_2392_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2392_word_address_0;
      ptr_deref_2392_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2414_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2414_store_0_req_0;
      ptr_deref_2414_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2414_store_0_req_1;
      ptr_deref_2414_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2414_word_address_0;
      data_in <= ptr_deref_2414_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2158_inst RPIPE_Block2_start_2161_inst RPIPE_Block2_start_2164_inst RPIPE_Block2_start_2167_inst RPIPE_Block2_start_2170_inst RPIPE_Block2_start_2173_inst RPIPE_Block2_start_2176_inst RPIPE_Block2_start_2179_inst RPIPE_Block2_start_2182_inst RPIPE_Block2_start_2185_inst RPIPE_Block2_start_2198_inst RPIPE_Block2_start_2210_inst RPIPE_Block2_start_2213_inst RPIPE_Block2_start_2216_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block2_start_2158_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2161_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2164_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2167_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2170_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2173_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2176_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2179_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2182_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2185_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2198_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2210_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2213_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2216_inst_req_0;
      RPIPE_Block2_start_2158_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2161_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2164_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2167_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2170_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2173_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2176_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2179_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2182_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2185_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2198_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2210_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2213_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2216_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block2_start_2158_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2161_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2164_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2167_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2170_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2173_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2176_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2179_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2182_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2185_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2198_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2210_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2213_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2216_inst_req_1;
      RPIPE_Block2_start_2158_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2161_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2164_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2167_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2170_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2173_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2176_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2179_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2182_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2185_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2198_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2210_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2213_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2216_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2159 <= data_out(223 downto 208);
      call1_2162 <= data_out(207 downto 192);
      call3_2165 <= data_out(191 downto 176);
      call5_2168 <= data_out(175 downto 160);
      call7_2171 <= data_out(159 downto 144);
      call9_2174 <= data_out(143 downto 128);
      call11_2177 <= data_out(127 downto 112);
      call13_2180 <= data_out(111 downto 96);
      call14_2183 <= data_out(95 downto 80);
      call15_2186 <= data_out(79 downto 64);
      call16_2199 <= data_out(63 downto 48);
      call18_2211 <= data_out(47 downto 32);
      call20_2214 <= data_out(31 downto 16);
      call22_2217 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2519_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2519_inst_req_0;
      WPIPE_Block2_done_2519_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2519_inst_req_1;
      WPIPE_Block2_done_2519_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2521_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6661_start: Boolean;
  signal convTransposeD_CP_6661_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2705_inst_ack_1 : boolean;
  signal addr_of_2773_final_reg_ack_0 : boolean;
  signal type_cast_2705_inst_req_1 : boolean;
  signal type_cast_2743_inst_req_0 : boolean;
  signal type_cast_2743_inst_ack_0 : boolean;
  signal addr_of_2750_final_reg_req_1 : boolean;
  signal ptr_deref_2754_load_0_req_1 : boolean;
  signal addr_of_2750_final_reg_ack_1 : boolean;
  signal ptr_deref_2754_load_0_ack_1 : boolean;
  signal addr_of_2773_final_reg_req_1 : boolean;
  signal type_cast_2713_inst_req_0 : boolean;
  signal type_cast_2743_inst_req_1 : boolean;
  signal type_cast_2743_inst_ack_1 : boolean;
  signal type_cast_2713_inst_ack_0 : boolean;
  signal addr_of_2773_final_reg_ack_1 : boolean;
  signal type_cast_2713_inst_req_1 : boolean;
  signal array_obj_ref_2749_index_offset_req_0 : boolean;
  signal array_obj_ref_2749_index_offset_ack_0 : boolean;
  signal type_cast_2713_inst_ack_1 : boolean;
  signal type_cast_2781_inst_req_1 : boolean;
  signal type_cast_2822_inst_ack_0 : boolean;
  signal type_cast_2781_inst_ack_1 : boolean;
  signal type_cast_2781_inst_req_0 : boolean;
  signal ptr_deref_2776_store_0_req_0 : boolean;
  signal ptr_deref_2776_store_0_req_1 : boolean;
  signal ptr_deref_2776_store_0_ack_1 : boolean;
  signal ptr_deref_2776_store_0_ack_0 : boolean;
  signal type_cast_2709_inst_req_0 : boolean;
  signal if_stmt_2794_branch_ack_1 : boolean;
  signal type_cast_2781_inst_ack_0 : boolean;
  signal type_cast_2822_inst_req_0 : boolean;
  signal if_stmt_2794_branch_ack_0 : boolean;
  signal if_stmt_2794_branch_req_0 : boolean;
  signal array_obj_ref_2772_index_offset_req_0 : boolean;
  signal RPIPE_Block3_start_2530_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2530_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2530_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2530_inst_ack_1 : boolean;
  signal type_cast_2709_inst_ack_1 : boolean;
  signal type_cast_2709_inst_req_1 : boolean;
  signal type_cast_2709_inst_ack_0 : boolean;
  signal addr_of_2750_final_reg_ack_0 : boolean;
  signal addr_of_2750_final_reg_req_0 : boolean;
  signal RPIPE_Block3_start_2533_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2533_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2533_inst_req_1 : boolean;
  signal ptr_deref_2754_load_0_ack_0 : boolean;
  signal RPIPE_Block3_start_2533_inst_ack_1 : boolean;
  signal addr_of_2773_final_reg_req_0 : boolean;
  signal RPIPE_Block3_start_2536_inst_req_0 : boolean;
  signal ptr_deref_2754_load_0_req_0 : boolean;
  signal RPIPE_Block3_start_2536_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2536_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2536_inst_ack_1 : boolean;
  signal array_obj_ref_2772_index_offset_ack_1 : boolean;
  signal RPIPE_Block3_start_2539_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2539_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2539_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2539_inst_ack_1 : boolean;
  signal array_obj_ref_2772_index_offset_req_1 : boolean;
  signal array_obj_ref_2772_index_offset_ack_0 : boolean;
  signal array_obj_ref_2749_index_offset_ack_1 : boolean;
  signal array_obj_ref_2749_index_offset_req_1 : boolean;
  signal RPIPE_Block3_start_2542_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2542_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2542_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2542_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2545_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2545_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2545_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2545_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2548_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2548_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2548_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2548_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2551_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2551_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2551_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2551_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2554_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2554_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2554_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2554_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2557_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2557_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2557_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2557_inst_ack_1 : boolean;
  signal type_cast_2561_inst_req_0 : boolean;
  signal type_cast_2561_inst_ack_0 : boolean;
  signal type_cast_2561_inst_req_1 : boolean;
  signal type_cast_2561_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2570_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2570_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2570_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2570_inst_ack_1 : boolean;
  signal type_cast_2574_inst_req_0 : boolean;
  signal type_cast_2574_inst_ack_0 : boolean;
  signal type_cast_2574_inst_req_1 : boolean;
  signal type_cast_2574_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2582_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2582_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2582_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2582_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2585_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2585_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2585_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2585_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2588_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2588_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2588_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2588_inst_ack_1 : boolean;
  signal type_cast_2632_inst_req_0 : boolean;
  signal type_cast_2632_inst_ack_0 : boolean;
  signal type_cast_2632_inst_req_1 : boolean;
  signal type_cast_2632_inst_ack_1 : boolean;
  signal type_cast_2636_inst_req_0 : boolean;
  signal type_cast_2636_inst_ack_0 : boolean;
  signal type_cast_2636_inst_req_1 : boolean;
  signal type_cast_2636_inst_ack_1 : boolean;
  signal type_cast_2640_inst_req_0 : boolean;
  signal type_cast_2640_inst_ack_0 : boolean;
  signal type_cast_2640_inst_req_1 : boolean;
  signal type_cast_2640_inst_ack_1 : boolean;
  signal type_cast_2705_inst_req_0 : boolean;
  signal type_cast_2705_inst_ack_0 : boolean;
  signal type_cast_2822_inst_req_1 : boolean;
  signal type_cast_2822_inst_ack_1 : boolean;
  signal if_stmt_2841_branch_req_0 : boolean;
  signal if_stmt_2841_branch_ack_1 : boolean;
  signal if_stmt_2841_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2877_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2877_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2877_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2877_inst_ack_1 : boolean;
  signal phi_stmt_2644_req_0 : boolean;
  signal phi_stmt_2651_req_0 : boolean;
  signal phi_stmt_2658_req_0 : boolean;
  signal type_cast_2668_inst_req_0 : boolean;
  signal type_cast_2668_inst_ack_0 : boolean;
  signal type_cast_2668_inst_req_1 : boolean;
  signal type_cast_2668_inst_ack_1 : boolean;
  signal phi_stmt_2665_req_0 : boolean;
  signal type_cast_2650_inst_req_0 : boolean;
  signal type_cast_2650_inst_ack_0 : boolean;
  signal type_cast_2650_inst_req_1 : boolean;
  signal type_cast_2650_inst_ack_1 : boolean;
  signal phi_stmt_2644_req_1 : boolean;
  signal type_cast_2657_inst_req_0 : boolean;
  signal type_cast_2657_inst_ack_0 : boolean;
  signal type_cast_2657_inst_req_1 : boolean;
  signal type_cast_2657_inst_ack_1 : boolean;
  signal phi_stmt_2651_req_1 : boolean;
  signal type_cast_2664_inst_req_0 : boolean;
  signal type_cast_2664_inst_ack_0 : boolean;
  signal type_cast_2664_inst_req_1 : boolean;
  signal type_cast_2664_inst_ack_1 : boolean;
  signal phi_stmt_2658_req_1 : boolean;
  signal type_cast_2670_inst_req_0 : boolean;
  signal type_cast_2670_inst_ack_0 : boolean;
  signal type_cast_2670_inst_req_1 : boolean;
  signal type_cast_2670_inst_ack_1 : boolean;
  signal phi_stmt_2665_req_1 : boolean;
  signal phi_stmt_2644_ack_0 : boolean;
  signal phi_stmt_2651_ack_0 : boolean;
  signal phi_stmt_2658_ack_0 : boolean;
  signal phi_stmt_2665_ack_0 : boolean;
  signal phi_stmt_2848_req_1 : boolean;
  signal type_cast_2860_inst_req_0 : boolean;
  signal type_cast_2860_inst_ack_0 : boolean;
  signal type_cast_2860_inst_req_1 : boolean;
  signal type_cast_2860_inst_ack_1 : boolean;
  signal phi_stmt_2855_req_1 : boolean;
  signal type_cast_2866_inst_req_0 : boolean;
  signal type_cast_2866_inst_ack_0 : boolean;
  signal type_cast_2866_inst_req_1 : boolean;
  signal type_cast_2866_inst_ack_1 : boolean;
  signal phi_stmt_2861_req_1 : boolean;
  signal type_cast_2851_inst_req_0 : boolean;
  signal type_cast_2851_inst_ack_0 : boolean;
  signal type_cast_2851_inst_req_1 : boolean;
  signal type_cast_2851_inst_ack_1 : boolean;
  signal phi_stmt_2848_req_0 : boolean;
  signal type_cast_2858_inst_req_0 : boolean;
  signal type_cast_2858_inst_ack_0 : boolean;
  signal type_cast_2858_inst_req_1 : boolean;
  signal type_cast_2858_inst_ack_1 : boolean;
  signal phi_stmt_2855_req_0 : boolean;
  signal type_cast_2864_inst_req_0 : boolean;
  signal type_cast_2864_inst_ack_0 : boolean;
  signal type_cast_2864_inst_req_1 : boolean;
  signal type_cast_2864_inst_ack_1 : boolean;
  signal phi_stmt_2861_req_0 : boolean;
  signal phi_stmt_2848_ack_0 : boolean;
  signal phi_stmt_2855_ack_0 : boolean;
  signal phi_stmt_2861_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6661_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6661_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6661_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6661_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6661: Block -- control-path 
    signal convTransposeD_CP_6661_elements: BooleanArray(123 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6661_elements(0) <= convTransposeD_CP_6661_start;
    convTransposeD_CP_6661_symbol <= convTransposeD_CP_6661_elements(74);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2528/$entry
      -- CP-element group 0: 	 branch_block_stmt_2528/branch_block_stmt_2528__entry__
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/$entry
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_Update/cr
      -- 
    rr_6709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(0), ack => RPIPE_Block3_start_2530_inst_req_0); -- 
    cr_6854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(0), ack => type_cast_2561_inst_req_1); -- 
    cr_6882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(0), ack => type_cast_2574_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	123 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	82 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2528/merge_stmt_2847__exit__
      -- CP-element group 1: 	 branch_block_stmt_2528/assign_stmt_2873__entry__
      -- CP-element group 1: 	 branch_block_stmt_2528/assign_stmt_2873__exit__
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2528/assign_stmt_2873/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/assign_stmt_2873/$exit
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/SplitProtocol/Update/cr
      -- 
    rr_7382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(1), ack => type_cast_2650_inst_req_0); -- 
    cr_7387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(1), ack => type_cast_2650_inst_req_1); -- 
    rr_7405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(1), ack => type_cast_2657_inst_req_0); -- 
    cr_7410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(1), ack => type_cast_2657_inst_req_1); -- 
    rr_7428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(1), ack => type_cast_2664_inst_req_0); -- 
    cr_7433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(1), ack => type_cast_2664_inst_req_1); -- 
    rr_7451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(1), ack => type_cast_2670_inst_req_0); -- 
    cr_7456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(1), ack => type_cast_2670_inst_req_1); -- 
    convTransposeD_CP_6661_elements(1) <= convTransposeD_CP_6661_elements(123);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_Update/cr
      -- 
    ra_6710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2530_inst_ack_0, ack => convTransposeD_CP_6661_elements(2)); -- 
    cr_6714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(2), ack => RPIPE_Block3_start_2530_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2530_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_Sample/rr
      -- 
    ca_6715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2530_inst_ack_1, ack => convTransposeD_CP_6661_elements(3)); -- 
    rr_6723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(3), ack => RPIPE_Block3_start_2533_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_Update/cr
      -- 
    ra_6724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2533_inst_ack_0, ack => convTransposeD_CP_6661_elements(4)); -- 
    cr_6728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(4), ack => RPIPE_Block3_start_2533_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2533_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_Sample/rr
      -- 
    ca_6729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2533_inst_ack_1, ack => convTransposeD_CP_6661_elements(5)); -- 
    rr_6737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(5), ack => RPIPE_Block3_start_2536_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_Update/cr
      -- 
    ra_6738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2536_inst_ack_0, ack => convTransposeD_CP_6661_elements(6)); -- 
    cr_6742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(6), ack => RPIPE_Block3_start_2536_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2536_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_Sample/rr
      -- 
    ca_6743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2536_inst_ack_1, ack => convTransposeD_CP_6661_elements(7)); -- 
    rr_6751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(7), ack => RPIPE_Block3_start_2539_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_Update/cr
      -- 
    ra_6752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2539_inst_ack_0, ack => convTransposeD_CP_6661_elements(8)); -- 
    cr_6756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(8), ack => RPIPE_Block3_start_2539_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2539_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_Sample/rr
      -- 
    ca_6757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2539_inst_ack_1, ack => convTransposeD_CP_6661_elements(9)); -- 
    rr_6765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(9), ack => RPIPE_Block3_start_2542_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_Update/cr
      -- 
    ra_6766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2542_inst_ack_0, ack => convTransposeD_CP_6661_elements(10)); -- 
    cr_6770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(10), ack => RPIPE_Block3_start_2542_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2542_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_Sample/rr
      -- 
    ca_6771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2542_inst_ack_1, ack => convTransposeD_CP_6661_elements(11)); -- 
    rr_6779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(11), ack => RPIPE_Block3_start_2545_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_Update/cr
      -- 
    ra_6780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2545_inst_ack_0, ack => convTransposeD_CP_6661_elements(12)); -- 
    cr_6784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(12), ack => RPIPE_Block3_start_2545_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2545_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_Sample/rr
      -- 
    ca_6785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2545_inst_ack_1, ack => convTransposeD_CP_6661_elements(13)); -- 
    rr_6793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(13), ack => RPIPE_Block3_start_2548_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_Update/cr
      -- 
    ra_6794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2548_inst_ack_0, ack => convTransposeD_CP_6661_elements(14)); -- 
    cr_6798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(14), ack => RPIPE_Block3_start_2548_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2548_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_Sample/rr
      -- 
    ca_6799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2548_inst_ack_1, ack => convTransposeD_CP_6661_elements(15)); -- 
    rr_6807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(15), ack => RPIPE_Block3_start_2551_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_Update/cr
      -- 
    ra_6808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2551_inst_ack_0, ack => convTransposeD_CP_6661_elements(16)); -- 
    cr_6812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(16), ack => RPIPE_Block3_start_2551_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2551_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_Sample/rr
      -- 
    ca_6813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2551_inst_ack_1, ack => convTransposeD_CP_6661_elements(17)); -- 
    rr_6821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(17), ack => RPIPE_Block3_start_2554_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_Update/cr
      -- 
    ra_6822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2554_inst_ack_0, ack => convTransposeD_CP_6661_elements(18)); -- 
    cr_6826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(18), ack => RPIPE_Block3_start_2554_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2554_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_Sample/rr
      -- 
    ca_6827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2554_inst_ack_1, ack => convTransposeD_CP_6661_elements(19)); -- 
    rr_6835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(19), ack => RPIPE_Block3_start_2557_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_Update/cr
      -- 
    ra_6836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2557_inst_ack_0, ack => convTransposeD_CP_6661_elements(20)); -- 
    cr_6840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(20), ack => RPIPE_Block3_start_2557_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2557_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_Sample/rr
      -- 
    ca_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2557_inst_ack_1, ack => convTransposeD_CP_6661_elements(21)); -- 
    rr_6849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(21), ack => type_cast_2561_inst_req_0); -- 
    rr_6863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(21), ack => RPIPE_Block3_start_2570_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_Sample/ra
      -- 
    ra_6850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2561_inst_ack_0, ack => convTransposeD_CP_6661_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2561_Update/ca
      -- 
    ca_6855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2561_inst_ack_1, ack => convTransposeD_CP_6661_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_Update/cr
      -- 
    ra_6864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2570_inst_ack_0, ack => convTransposeD_CP_6661_elements(24)); -- 
    cr_6868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(24), ack => RPIPE_Block3_start_2570_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2570_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_Sample/rr
      -- 
    ca_6869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2570_inst_ack_1, ack => convTransposeD_CP_6661_elements(25)); -- 
    rr_6877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(25), ack => type_cast_2574_inst_req_0); -- 
    rr_6891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(25), ack => RPIPE_Block3_start_2582_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_Sample/ra
      -- 
    ra_6878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2574_inst_ack_0, ack => convTransposeD_CP_6661_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/type_cast_2574_Update/ca
      -- 
    ca_6883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2574_inst_ack_1, ack => convTransposeD_CP_6661_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_Update/cr
      -- 
    ra_6892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2582_inst_ack_0, ack => convTransposeD_CP_6661_elements(28)); -- 
    cr_6896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(28), ack => RPIPE_Block3_start_2582_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2582_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_Sample/rr
      -- 
    ca_6897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2582_inst_ack_1, ack => convTransposeD_CP_6661_elements(29)); -- 
    rr_6905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(29), ack => RPIPE_Block3_start_2585_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_Update/cr
      -- 
    ra_6906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2585_inst_ack_0, ack => convTransposeD_CP_6661_elements(30)); -- 
    cr_6910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(30), ack => RPIPE_Block3_start_2585_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2585_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_Sample/rr
      -- 
    ca_6911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2585_inst_ack_1, ack => convTransposeD_CP_6661_elements(31)); -- 
    rr_6919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(31), ack => RPIPE_Block3_start_2588_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_Update/cr
      -- 
    ra_6920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2588_inst_ack_0, ack => convTransposeD_CP_6661_elements(32)); -- 
    cr_6924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(32), ack => RPIPE_Block3_start_2588_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/RPIPE_Block3_start_2588_Update/ca
      -- 
    ca_6925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2588_inst_ack_1, ack => convTransposeD_CP_6661_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589__exit__
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641__entry__
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2531_to_assign_stmt_2589/$exit
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/$entry
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_Update/cr
      -- 
    rr_6936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(34), ack => type_cast_2632_inst_req_0); -- 
    cr_6941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(34), ack => type_cast_2632_inst_req_1); -- 
    rr_6950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(34), ack => type_cast_2636_inst_req_0); -- 
    cr_6955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(34), ack => type_cast_2636_inst_req_1); -- 
    rr_6964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(34), ack => type_cast_2640_inst_req_0); -- 
    cr_6969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(34), ack => type_cast_2640_inst_req_1); -- 
    convTransposeD_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(23) & convTransposeD_CP_6661_elements(27) & convTransposeD_CP_6661_elements(33);
      gj_convTransposeD_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_Sample/ra
      -- 
    ra_6937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2632_inst_ack_0, ack => convTransposeD_CP_6661_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	41 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2632_Update/ca
      -- 
    ca_6942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2632_inst_ack_1, ack => convTransposeD_CP_6661_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_Sample/ra
      -- 
    ra_6951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2636_inst_ack_0, ack => convTransposeD_CP_6661_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2636_Update/ca
      -- 
    ca_6956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2636_inst_ack_1, ack => convTransposeD_CP_6661_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_Sample/ra
      -- 
    ra_6965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2640_inst_ack_0, ack => convTransposeD_CP_6661_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/type_cast_2640_Update/ca
      -- 
    ca_6970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2640_inst_ack_1, ack => convTransposeD_CP_6661_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	36 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	75 
    -- CP-element group 41: 	76 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	78 
    -- CP-element group 41: 	79 
    -- CP-element group 41:  members (18) 
      -- CP-element group 41: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641__exit__
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody
      -- CP-element group 41: 	 branch_block_stmt_2528/assign_stmt_2596_to_assign_stmt_2641/$exit
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2644/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2651/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2658/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/SplitProtocol/Update/cr
      -- 
    rr_7356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(41), ack => type_cast_2668_inst_req_0); -- 
    cr_7361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(41), ack => type_cast_2668_inst_req_1); -- 
    convTransposeD_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(36) & convTransposeD_CP_6661_elements(38) & convTransposeD_CP_6661_elements(40);
      gj_convTransposeD_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	100 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_Sample/ra
      -- 
    ra_6982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2705_inst_ack_0, ack => convTransposeD_CP_6661_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	100 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_Update/$exit
      -- 
    ca_6987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2705_inst_ack_1, ack => convTransposeD_CP_6661_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	100 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_Sample/ra
      -- 
    ra_6996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_0, ack => convTransposeD_CP_6661_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	100 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	56 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_Update/$exit
      -- 
    ca_7001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_1, ack => convTransposeD_CP_6661_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	100 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_Sample/ra
      -- 
    ra_7010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2713_inst_ack_0, ack => convTransposeD_CP_6661_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	100 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_Update/ca
      -- 
    ca_7015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2713_inst_ack_1, ack => convTransposeD_CP_6661_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	100 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_sample_completed_
      -- 
    ra_7024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2743_inst_ack_0, ack => convTransposeD_CP_6661_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	100 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_final_index_sum_regn_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_update_completed_
      -- 
    ca_7029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2743_inst_ack_1, ack => convTransposeD_CP_6661_elements(49)); -- 
    req_7054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(49), ack => array_obj_ref_2749_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	66 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_final_index_sum_regn_sample_complete
      -- CP-element group 50: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_final_index_sum_regn_Sample/ack
      -- 
    ack_7055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2749_index_offset_ack_0, ack => convTransposeD_CP_6661_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	100 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_request/req
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_base_plus_offset/sum_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_final_index_sum_regn_Update/$exit
      -- 
    ack_7060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2749_index_offset_ack_1, ack => convTransposeD_CP_6661_elements(51)); -- 
    req_7069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(51), ack => addr_of_2750_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_request/ack
      -- CP-element group 52: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_request/$exit
      -- 
    ack_7070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2750_final_reg_ack_0, ack => convTransposeD_CP_6661_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	100 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (24) 
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Sample/word_access_start/word_0/rr
      -- CP-element group 53: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Sample/word_access_start/word_0/$entry
      -- 
    ack_7075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2750_final_reg_ack_1, ack => convTransposeD_CP_6661_elements(53)); -- 
    rr_7108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(53), ack => ptr_deref_2754_load_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Sample/word_access_start/word_0/ra
      -- CP-element group 54: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Sample/word_access_start/$exit
      -- 
    ra_7109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2754_load_0_ack_0, ack => convTransposeD_CP_6661_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	100 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/ptr_deref_2754_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/ptr_deref_2754_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/ptr_deref_2754_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/ptr_deref_2754_Merge/merge_ack
      -- CP-element group 55: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/$exit
      -- 
    ca_7120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2754_load_0_ack_1, ack => convTransposeD_CP_6661_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	45 
    -- CP-element group 56: 	47 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (13) 
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_final_index_sum_regn_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_index_resize_1/$exit
      -- 
    req_7150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(56), ack => array_obj_ref_2772_index_offset_req_0); -- 
    convTransposeD_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(43) & convTransposeD_CP_6661_elements(45) & convTransposeD_CP_6661_elements(47);
      gj_convTransposeD_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_final_index_sum_regn_Sample/ack
      -- 
    ack_7151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2772_index_offset_ack_0, ack => convTransposeD_CP_6661_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	100 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_request/req
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_final_index_sum_regn_Update/$exit
      -- 
    ack_7156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2772_index_offset_ack_1, ack => convTransposeD_CP_6661_elements(58)); -- 
    req_7165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(58), ack => addr_of_2773_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_request/ack
      -- CP-element group 59: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_request/$exit
      -- 
    ack_7166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2773_final_reg_ack_0, ack => convTransposeD_CP_6661_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	100 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (19) 
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_word_addrgen/root_register_ack
      -- 
    ack_7171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2773_final_reg_ack_1, ack => convTransposeD_CP_6661_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/ptr_deref_2776_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/ptr_deref_2776_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/word_access_start/word_0/rr
      -- CP-element group 61: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/ptr_deref_2776_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/ptr_deref_2776_Split/$entry
      -- 
    rr_7209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(61), ack => ptr_deref_2776_store_0_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(55) & convTransposeD_CP_6661_elements(60);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Sample/word_access_start/word_0/ra
      -- 
    ra_7210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2776_store_0_ack_0, ack => convTransposeD_CP_6661_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	100 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Update/word_access_complete/word_0/ca
      -- 
    ca_7221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2776_store_0_ack_1, ack => convTransposeD_CP_6661_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	100 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_Sample/ra
      -- 
    ra_7230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2781_inst_ack_0, ack => convTransposeD_CP_6661_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	100 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_Update/ca
      -- CP-element group 65: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_update_completed_
      -- 
    ca_7235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2781_inst_ack_1, ack => convTransposeD_CP_6661_elements(65)); -- 
    -- CP-element group 66:  branch  join  transition  place  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	50 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	63 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (10) 
      -- CP-element group 66: 	 branch_block_stmt_2528/if_stmt_2794__entry__
      -- CP-element group 66: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793__exit__
      -- CP-element group 66: 	 branch_block_stmt_2528/R_cmp_2795_place
      -- CP-element group 66: 	 branch_block_stmt_2528/if_stmt_2794_else_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2528/if_stmt_2794_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2528/if_stmt_2794_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2528/if_stmt_2794_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2528/if_stmt_2794_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2528/if_stmt_2794_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/$exit
      -- 
    branch_req_7243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(66), ack => if_stmt_2794_branch_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(50) & convTransposeD_CP_6661_elements(57) & convTransposeD_CP_6661_elements(63) & convTransposeD_CP_6661_elements(65);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	109 
    -- CP-element group 67: 	110 
    -- CP-element group 67: 	112 
    -- CP-element group 67: 	113 
    -- CP-element group 67: 	115 
    -- CP-element group 67: 	116 
    -- CP-element group 67:  members (40) 
      -- CP-element group 67: 	 branch_block_stmt_2528/whilex_xbody_ifx_xthen
      -- CP-element group 67: 	 branch_block_stmt_2528/merge_stmt_2800__exit__
      -- CP-element group 67: 	 branch_block_stmt_2528/assign_stmt_2806__entry__
      -- CP-element group 67: 	 branch_block_stmt_2528/assign_stmt_2806__exit__
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132
      -- CP-element group 67: 	 branch_block_stmt_2528/merge_stmt_2800_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2528/if_stmt_2794_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2528/assign_stmt_2806/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/assign_stmt_2806/$exit
      -- CP-element group 67: 	 branch_block_stmt_2528/if_stmt_2794_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2528/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2528/merge_stmt_2800_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/merge_stmt_2800_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2528/merge_stmt_2800_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2794_branch_ack_1, ack => convTransposeD_CP_6661_elements(67)); -- 
    rr_7566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(67), ack => type_cast_2851_inst_req_0); -- 
    cr_7571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(67), ack => type_cast_2851_inst_req_1); -- 
    rr_7589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(67), ack => type_cast_2858_inst_req_0); -- 
    cr_7594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(67), ack => type_cast_2858_inst_req_1); -- 
    rr_7612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(67), ack => type_cast_2864_inst_req_0); -- 
    cr_7617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(67), ack => type_cast_2864_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (18) 
      -- CP-element group 68: 	 branch_block_stmt_2528/whilex_xbody_ifx_xelse
      -- CP-element group 68: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840__entry__
      -- CP-element group 68: 	 branch_block_stmt_2528/merge_stmt_2808__exit__
      -- CP-element group 68: 	 branch_block_stmt_2528/merge_stmt_2808_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/$entry
      -- CP-element group 68: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_update_start_
      -- CP-element group 68: 	 branch_block_stmt_2528/if_stmt_2794_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2528/if_stmt_2794_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2528/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2528/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_2528/merge_stmt_2808_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_2528/merge_stmt_2808_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_2528/merge_stmt_2808_PhiAck/dummy
      -- 
    else_choice_transition_7252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2794_branch_ack_0, ack => convTransposeD_CP_6661_elements(68)); -- 
    rr_7268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(68), ack => type_cast_2822_inst_req_0); -- 
    cr_7273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(68), ack => type_cast_2822_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_Sample/$exit
      -- 
    ra_7269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2822_inst_ack_0, ack => convTransposeD_CP_6661_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2528/R_cmp121_2842_place
      -- CP-element group 70: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840__exit__
      -- CP-element group 70: 	 branch_block_stmt_2528/if_stmt_2841__entry__
      -- CP-element group 70: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/$exit
      -- CP-element group 70: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2528/assign_stmt_2814_to_assign_stmt_2840/type_cast_2822_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2528/if_stmt_2841_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2528/if_stmt_2841_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2528/if_stmt_2841_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2528/if_stmt_2841_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2528/if_stmt_2841_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2528/if_stmt_2841_else_link/$entry
      -- 
    ca_7274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2822_inst_ack_1, ack => convTransposeD_CP_6661_elements(70)); -- 
    branch_req_7282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(70), ack => if_stmt_2841_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2528/ifx_xelse_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2528/merge_stmt_2875_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2528/merge_stmt_2875__exit__
      -- CP-element group 71: 	 branch_block_stmt_2528/assign_stmt_2880__entry__
      -- CP-element group 71: 	 branch_block_stmt_2528/if_stmt_2841_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2528/if_stmt_2841_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2528/assign_stmt_2880/$entry
      -- CP-element group 71: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2528/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2528/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2528/merge_stmt_2875_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2528/merge_stmt_2875_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2528/merge_stmt_2875_PhiAck/dummy
      -- 
    if_choice_transition_7287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2841_branch_ack_1, ack => convTransposeD_CP_6661_elements(71)); -- 
    req_7307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(71), ack => WPIPE_Block3_done_2877_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	101 
    -- CP-element group 72: 	102 
    -- CP-element group 72: 	103 
    -- CP-element group 72: 	105 
    -- CP-element group 72: 	106 
    -- CP-element group 72:  members (22) 
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/if_stmt_2841_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2528/if_stmt_2841_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2848/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2841_branch_ack_0, ack => convTransposeD_CP_6661_elements(72)); -- 
    rr_7517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(72), ack => type_cast_2860_inst_req_0); -- 
    cr_7522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(72), ack => type_cast_2860_inst_req_1); -- 
    rr_7540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(72), ack => type_cast_2866_inst_req_0); -- 
    cr_7545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(72), ack => type_cast_2866_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_Update/req
      -- 
    ack_7308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2877_inst_ack_0, ack => convTransposeD_CP_6661_elements(73)); -- 
    req_7312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(73), ack => WPIPE_Block3_done_2877_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 branch_block_stmt_2528/merge_stmt_2882_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2528/branch_block_stmt_2528__exit__
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2528/$exit
      -- CP-element group 74: 	 branch_block_stmt_2528/assign_stmt_2880__exit__
      -- CP-element group 74: 	 branch_block_stmt_2528/return__
      -- CP-element group 74: 	 branch_block_stmt_2528/merge_stmt_2882__exit__
      -- CP-element group 74: 	 branch_block_stmt_2528/assign_stmt_2880/$exit
      -- CP-element group 74: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2528/assign_stmt_2880/WPIPE_Block3_done_2877_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2528/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2528/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2528/merge_stmt_2882_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2528/merge_stmt_2882_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2528/merge_stmt_2882_PhiAck/dummy
      -- 
    ack_7313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2877_inst_ack_1, ack => convTransposeD_CP_6661_elements(74)); -- 
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	81 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2644/$exit
      -- CP-element group 75: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2648_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_req
      -- 
    phi_stmt_2644_req_7324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2644_req_7324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(75), ack => phi_stmt_2644_req_0); -- 
    -- Element group convTransposeD_CP_6661_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeD_CP_6661_elements(41), ack => convTransposeD_CP_6661_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  output  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	41 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	81 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2651/$exit
      -- CP-element group 76: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2655_konst_delay_trans
      -- CP-element group 76: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_req
      -- 
    phi_stmt_2651_req_7332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2651_req_7332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(76), ack => phi_stmt_2651_req_0); -- 
    -- Element group convTransposeD_CP_6661_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => convTransposeD_CP_6661_elements(41), ack => convTransposeD_CP_6661_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	41 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2658/$exit
      -- CP-element group 77: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2662_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_req
      -- 
    phi_stmt_2658_req_7340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2658_req_7340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(77), ack => phi_stmt_2658_req_0); -- 
    -- Element group convTransposeD_CP_6661_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeD_CP_6661_elements(41), ack => convTransposeD_CP_6661_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	41 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/SplitProtocol/Sample/ra
      -- 
    ra_7357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2668_inst_ack_0, ack => convTransposeD_CP_6661_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	41 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/SplitProtocol/Update/ca
      -- 
    ca_7362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2668_inst_ack_1, ack => convTransposeD_CP_6661_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/$exit
      -- CP-element group 80: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/$exit
      -- CP-element group 80: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2668/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_req
      -- 
    phi_stmt_2665_req_7363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2665_req_7363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(80), ack => phi_stmt_2665_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(78) & convTransposeD_CP_6661_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: 	76 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	95 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2528/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(75) & convTransposeD_CP_6661_elements(76) & convTransposeD_CP_6661_elements(77) & convTransposeD_CP_6661_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	1 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/SplitProtocol/Sample/ra
      -- 
    ra_7383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2650_inst_ack_0, ack => convTransposeD_CP_6661_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/SplitProtocol/Update/ca
      -- 
    ca_7388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2650_inst_ack_1, ack => convTransposeD_CP_6661_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	94 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/$exit
      -- CP-element group 84: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/$exit
      -- CP-element group 84: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_sources/type_cast_2650/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2644/phi_stmt_2644_req
      -- 
    phi_stmt_2644_req_7389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2644_req_7389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(84), ack => phi_stmt_2644_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(82) & convTransposeD_CP_6661_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/SplitProtocol/Sample/ra
      -- 
    ra_7406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2657_inst_ack_0, ack => convTransposeD_CP_6661_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/SplitProtocol/Update/ca
      -- 
    ca_7411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2657_inst_ack_1, ack => convTransposeD_CP_6661_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	94 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/$exit
      -- CP-element group 87: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/$exit
      -- CP-element group 87: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_sources/type_cast_2657/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2651/phi_stmt_2651_req
      -- 
    phi_stmt_2651_req_7412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2651_req_7412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(87), ack => phi_stmt_2651_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(85) & convTransposeD_CP_6661_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/SplitProtocol/Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/SplitProtocol/Sample/ra
      -- 
    ra_7429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2664_inst_ack_0, ack => convTransposeD_CP_6661_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/SplitProtocol/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/SplitProtocol/Update/ca
      -- 
    ca_7434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2664_inst_ack_1, ack => convTransposeD_CP_6661_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/$exit
      -- CP-element group 90: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/$exit
      -- CP-element group 90: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_sources/type_cast_2664/SplitProtocol/$exit
      -- CP-element group 90: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2658/phi_stmt_2658_req
      -- 
    phi_stmt_2658_req_7435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2658_req_7435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(90), ack => phi_stmt_2658_req_1); -- 
    convTransposeD_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(88) & convTransposeD_CP_6661_elements(89);
      gj_convTransposeD_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/SplitProtocol/Sample/ra
      -- 
    ra_7452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2670_inst_ack_0, ack => convTransposeD_CP_6661_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/SplitProtocol/Update/ca
      -- 
    ca_7457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2670_inst_ack_1, ack => convTransposeD_CP_6661_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/$exit
      -- CP-element group 93: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/$exit
      -- CP-element group 93: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_sources/type_cast_2670/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2665/phi_stmt_2665_req
      -- 
    phi_stmt_2665_req_7458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2665_req_7458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(93), ack => phi_stmt_2665_req_1); -- 
    convTransposeD_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(91) & convTransposeD_CP_6661_elements(92);
      gj_convTransposeD_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	84 
    -- CP-element group 94: 	87 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2528/ifx_xend132_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(84) & convTransposeD_CP_6661_elements(87) & convTransposeD_CP_6661_elements(90) & convTransposeD_CP_6661_elements(93);
      gj_convTransposeD_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  merge  fork  transition  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	81 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	98 
    -- CP-element group 95: 	99 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2528/merge_stmt_2643_PhiReqMerge
      -- CP-element group 95: 	 branch_block_stmt_2528/merge_stmt_2643_PhiAck/$entry
      -- 
    convTransposeD_CP_6661_elements(95) <= OrReduce(convTransposeD_CP_6661_elements(81) & convTransposeD_CP_6661_elements(94));
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2528/merge_stmt_2643_PhiAck/phi_stmt_2644_ack
      -- 
    phi_stmt_2644_ack_7463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2644_ack_0, ack => convTransposeD_CP_6661_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2528/merge_stmt_2643_PhiAck/phi_stmt_2651_ack
      -- 
    phi_stmt_2651_ack_7464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2651_ack_0, ack => convTransposeD_CP_6661_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2528/merge_stmt_2643_PhiAck/phi_stmt_2658_ack
      -- 
    phi_stmt_2658_ack_7465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2658_ack_0, ack => convTransposeD_CP_6661_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	95 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2528/merge_stmt_2643_PhiAck/phi_stmt_2665_ack
      -- 
    phi_stmt_2665_ack_7466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2665_ack_0, ack => convTransposeD_CP_6661_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  place  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	97 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	42 
    -- CP-element group 100: 	43 
    -- CP-element group 100: 	44 
    -- CP-element group 100: 	45 
    -- CP-element group 100: 	46 
    -- CP-element group 100: 	47 
    -- CP-element group 100: 	48 
    -- CP-element group 100: 	49 
    -- CP-element group 100: 	51 
    -- CP-element group 100: 	53 
    -- CP-element group 100: 	55 
    -- CP-element group 100: 	58 
    -- CP-element group 100: 	60 
    -- CP-element group 100: 	63 
    -- CP-element group 100: 	64 
    -- CP-element group 100: 	65 
    -- CP-element group 100:  members (56) 
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2528/merge_stmt_2643__exit__
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793__entry__
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2773_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/addr_of_2750_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2776_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2781_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2713_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2709_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/ptr_deref_2754_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2743_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2772_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/array_obj_ref_2749_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2528/assign_stmt_2677_to_assign_stmt_2793/type_cast_2705_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2528/merge_stmt_2643_PhiAck/$exit
      -- 
    cr_6986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => type_cast_2705_inst_req_1); -- 
    rr_7023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => type_cast_2743_inst_req_0); -- 
    req_7074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => addr_of_2750_final_reg_req_1); -- 
    cr_7119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => ptr_deref_2754_load_0_req_1); -- 
    req_7170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => addr_of_2773_final_reg_req_1); -- 
    rr_7009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => type_cast_2713_inst_req_0); -- 
    cr_7028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => type_cast_2743_inst_req_1); -- 
    cr_7014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => type_cast_2713_inst_req_1); -- 
    cr_7234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => type_cast_2781_inst_req_1); -- 
    rr_7229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => type_cast_2781_inst_req_0); -- 
    cr_7220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => ptr_deref_2776_store_0_req_1); -- 
    rr_6995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => type_cast_2709_inst_req_0); -- 
    cr_7000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => type_cast_2709_inst_req_1); -- 
    req_7155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => array_obj_ref_2772_index_offset_req_1); -- 
    req_7059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => array_obj_ref_2749_index_offset_req_1); -- 
    rr_6981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(100), ack => type_cast_2705_inst_req_0); -- 
    convTransposeD_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(96) & convTransposeD_CP_6661_elements(97) & convTransposeD_CP_6661_elements(98) & convTransposeD_CP_6661_elements(99);
      gj_convTransposeD_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  output  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	72 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2848/$exit
      -- CP-element group 101: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2854_konst_delay_trans
      -- CP-element group 101: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_req
      -- 
    phi_stmt_2848_req_7501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2848_req_7501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(101), ack => phi_stmt_2848_req_1); -- 
    -- Element group convTransposeD_CP_6661_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => convTransposeD_CP_6661_elements(72), ack => convTransposeD_CP_6661_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	72 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/SplitProtocol/Sample/ra
      -- 
    ra_7518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2860_inst_ack_0, ack => convTransposeD_CP_6661_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	72 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/SplitProtocol/Update/ca
      -- 
    ca_7523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2860_inst_ack_1, ack => convTransposeD_CP_6661_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/$exit
      -- CP-element group 104: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/$exit
      -- CP-element group 104: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2860/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_req
      -- 
    phi_stmt_2855_req_7524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2855_req_7524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(104), ack => phi_stmt_2855_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(102) & convTransposeD_CP_6661_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	72 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/SplitProtocol/Sample/ra
      -- 
    ra_7541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2866_inst_ack_0, ack => convTransposeD_CP_6661_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	72 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/SplitProtocol/Update/ca
      -- 
    ca_7546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2866_inst_ack_1, ack => convTransposeD_CP_6661_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/$exit
      -- CP-element group 107: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/$exit
      -- CP-element group 107: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2866/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_req
      -- 
    phi_stmt_2861_req_7547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2861_req_7547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(107), ack => phi_stmt_2861_req_1); -- 
    convTransposeD_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(105) & convTransposeD_CP_6661_elements(106);
      gj_convTransposeD_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2528/ifx_xelse_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(101) & convTransposeD_CP_6661_elements(104) & convTransposeD_CP_6661_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	67 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/SplitProtocol/Sample/ra
      -- 
    ra_7567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2851_inst_ack_0, ack => convTransposeD_CP_6661_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	67 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/SplitProtocol/Update/ca
      -- 
    ca_7572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2851_inst_ack_1, ack => convTransposeD_CP_6661_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	118 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/$exit
      -- CP-element group 111: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/$exit
      -- CP-element group 111: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_sources/type_cast_2851/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2848/phi_stmt_2848_req
      -- 
    phi_stmt_2848_req_7573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2848_req_7573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(111), ack => phi_stmt_2848_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(109) & convTransposeD_CP_6661_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/SplitProtocol/Sample/ra
      -- 
    ra_7590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2858_inst_ack_0, ack => convTransposeD_CP_6661_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	67 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/SplitProtocol/Update/ca
      -- 
    ca_7595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2858_inst_ack_1, ack => convTransposeD_CP_6661_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/$exit
      -- CP-element group 114: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/$exit
      -- CP-element group 114: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_sources/type_cast_2858/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2855/phi_stmt_2855_req
      -- 
    phi_stmt_2855_req_7596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2855_req_7596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(114), ack => phi_stmt_2855_req_0); -- 
    convTransposeD_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(112) & convTransposeD_CP_6661_elements(113);
      gj_convTransposeD_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	67 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/SplitProtocol/Sample/ra
      -- 
    ra_7613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2864_inst_ack_0, ack => convTransposeD_CP_6661_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	67 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/SplitProtocol/Update/ca
      -- 
    ca_7618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2864_inst_ack_1, ack => convTransposeD_CP_6661_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/$exit
      -- CP-element group 117: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/$exit
      -- CP-element group 117: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_sources/type_cast_2864/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2861/phi_stmt_2861_req
      -- 
    phi_stmt_2861_req_7619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2861_req_7619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6661_elements(117), ack => phi_stmt_2861_req_0); -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(115) & convTransposeD_CP_6661_elements(116);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	111 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2528/ifx_xthen_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(111) & convTransposeD_CP_6661_elements(114) & convTransposeD_CP_6661_elements(117);
      gj_convTransposeD_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2528/merge_stmt_2847_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_2528/merge_stmt_2847_PhiAck/$entry
      -- 
    convTransposeD_CP_6661_elements(119) <= OrReduce(convTransposeD_CP_6661_elements(108) & convTransposeD_CP_6661_elements(118));
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2528/merge_stmt_2847_PhiAck/phi_stmt_2848_ack
      -- 
    phi_stmt_2848_ack_7624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2848_ack_0, ack => convTransposeD_CP_6661_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_2528/merge_stmt_2847_PhiAck/phi_stmt_2855_ack
      -- 
    phi_stmt_2855_ack_7625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2855_ack_0, ack => convTransposeD_CP_6661_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2528/merge_stmt_2847_PhiAck/phi_stmt_2861_ack
      -- 
    phi_stmt_2861_ack_7626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2861_ack_0, ack => convTransposeD_CP_6661_elements(122)); -- 
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	120 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	1 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2528/merge_stmt_2847_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6661_elements(120) & convTransposeD_CP_6661_elements(121) & convTransposeD_CP_6661_elements(122);
      gj_convTransposeD_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6661_elements(123), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom91_2771_resized : std_logic_vector(13 downto 0);
    signal R_idxprom91_2771_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2748_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2748_scaled : std_logic_vector(13 downto 0);
    signal add103_2806 : std_logic_vector(15 downto 0);
    signal add32_2607 : std_logic_vector(15 downto 0);
    signal add50_2613 : std_logic_vector(15 downto 0);
    signal add63_2624 : std_logic_vector(15 downto 0);
    signal add82_2724 : std_logic_vector(63 downto 0);
    signal add84_2734 : std_logic_vector(63 downto 0);
    signal add96_2788 : std_logic_vector(31 downto 0);
    signal add_2580 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2682 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2749_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2749_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2749_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2749_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2749_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2749_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2772_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2772_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2772_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2772_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2772_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2772_root_address : std_logic_vector(13 downto 0);
    signal arrayidx87_2751 : std_logic_vector(31 downto 0);
    signal arrayidx92_2774 : std_logic_vector(31 downto 0);
    signal call11_2549 : std_logic_vector(15 downto 0);
    signal call13_2552 : std_logic_vector(15 downto 0);
    signal call14_2555 : std_logic_vector(15 downto 0);
    signal call15_2558 : std_logic_vector(15 downto 0);
    signal call16_2571 : std_logic_vector(15 downto 0);
    signal call18_2583 : std_logic_vector(15 downto 0);
    signal call1_2534 : std_logic_vector(15 downto 0);
    signal call20_2586 : std_logic_vector(15 downto 0);
    signal call22_2589 : std_logic_vector(15 downto 0);
    signal call3_2537 : std_logic_vector(15 downto 0);
    signal call5_2540 : std_logic_vector(15 downto 0);
    signal call7_2543 : std_logic_vector(15 downto 0);
    signal call9_2546 : std_logic_vector(15 downto 0);
    signal call_2531 : std_logic_vector(15 downto 0);
    signal cmp111_2819 : std_logic_vector(0 downto 0);
    signal cmp121_2840 : std_logic_vector(0 downto 0);
    signal cmp_2793 : std_logic_vector(0 downto 0);
    signal conv17_2575 : std_logic_vector(31 downto 0);
    signal conv70_2706 : std_logic_vector(63 downto 0);
    signal conv73_2633 : std_logic_vector(63 downto 0);
    signal conv75_2710 : std_logic_vector(63 downto 0);
    signal conv78_2637 : std_logic_vector(63 downto 0);
    signal conv80_2714 : std_logic_vector(63 downto 0);
    signal conv95_2782 : std_logic_vector(31 downto 0);
    signal conv99_2641 : std_logic_vector(31 downto 0);
    signal conv_2562 : std_logic_vector(31 downto 0);
    signal idxprom91_2767 : std_logic_vector(63 downto 0);
    signal idxprom_2744 : std_logic_vector(63 downto 0);
    signal inc115_2823 : std_logic_vector(15 downto 0);
    signal inc115x_xinput_dim0x_x2_2828 : std_logic_vector(15 downto 0);
    signal inc_2814 : std_logic_vector(15 downto 0);
    signal indvar_2644 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2873 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2861 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2665 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2855 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2658 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2835 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2848 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2651 : std_logic_vector(15 downto 0);
    signal mul59_2697 : std_logic_vector(15 downto 0);
    signal mul81_2719 : std_logic_vector(63 downto 0);
    signal mul83_2729 : std_logic_vector(63 downto 0);
    signal mul_2687 : std_logic_vector(15 downto 0);
    signal ptr_deref_2754_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2754_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2754_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2754_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2754_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2776_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2776_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2776_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2776_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2776_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2776_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2568 : std_logic_vector(31 downto 0);
    signal shr135_2596 : std_logic_vector(15 downto 0);
    signal shr31136_2602 : std_logic_vector(15 downto 0);
    signal shr86_2740 : std_logic_vector(31 downto 0);
    signal shr90_2761 : std_logic_vector(63 downto 0);
    signal sub53_2692 : std_logic_vector(15 downto 0);
    signal sub66_2629 : std_logic_vector(15 downto 0);
    signal sub67_2702 : std_logic_vector(15 downto 0);
    signal sub_2618 : std_logic_vector(15 downto 0);
    signal tmp1_2677 : std_logic_vector(31 downto 0);
    signal tmp88_2755 : std_logic_vector(63 downto 0);
    signal type_cast_2566_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2594_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2600_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2611_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2622_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2648_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2650_wire : std_logic_vector(31 downto 0);
    signal type_cast_2655_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2657_wire : std_logic_vector(15 downto 0);
    signal type_cast_2662_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2664_wire : std_logic_vector(15 downto 0);
    signal type_cast_2668_wire : std_logic_vector(15 downto 0);
    signal type_cast_2670_wire : std_logic_vector(15 downto 0);
    signal type_cast_2675_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2738_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2759_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2765_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2786_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2804_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2812_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2832_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2851_wire : std_logic_vector(15 downto 0);
    signal type_cast_2854_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2858_wire : std_logic_vector(15 downto 0);
    signal type_cast_2860_wire : std_logic_vector(15 downto 0);
    signal type_cast_2864_wire : std_logic_vector(15 downto 0);
    signal type_cast_2866_wire : std_logic_vector(15 downto 0);
    signal type_cast_2871_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2879_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2749_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2749_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2749_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2749_resized_base_address <= "00000000000000";
    array_obj_ref_2772_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2772_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2772_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2772_resized_base_address <= "00000000000000";
    ptr_deref_2754_word_offset_0 <= "00000000000000";
    ptr_deref_2776_word_offset_0 <= "00000000000000";
    type_cast_2566_wire_constant <= "00000000000000000000000000010000";
    type_cast_2594_wire_constant <= "0000000000000010";
    type_cast_2600_wire_constant <= "0000000000000001";
    type_cast_2611_wire_constant <= "1111111111111111";
    type_cast_2622_wire_constant <= "1111111111111111";
    type_cast_2648_wire_constant <= "00000000000000000000000000000000";
    type_cast_2655_wire_constant <= "0000000000000000";
    type_cast_2662_wire_constant <= "0000000000000000";
    type_cast_2675_wire_constant <= "00000000000000000000000000000100";
    type_cast_2738_wire_constant <= "00000000000000000000000000000010";
    type_cast_2759_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2765_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2786_wire_constant <= "00000000000000000000000000000100";
    type_cast_2804_wire_constant <= "0000000000000100";
    type_cast_2812_wire_constant <= "0000000000000001";
    type_cast_2832_wire_constant <= "0000000000000000";
    type_cast_2854_wire_constant <= "0000000000000000";
    type_cast_2871_wire_constant <= "00000000000000000000000000000001";
    type_cast_2879_wire_constant <= "0000000000000001";
    phi_stmt_2644: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2648_wire_constant & type_cast_2650_wire;
      req <= phi_stmt_2644_req_0 & phi_stmt_2644_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2644",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2644_ack_0,
          idata => idata,
          odata => indvar_2644,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2644
    phi_stmt_2651: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2655_wire_constant & type_cast_2657_wire;
      req <= phi_stmt_2651_req_0 & phi_stmt_2651_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2651",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2651_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2651,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2651
    phi_stmt_2658: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2662_wire_constant & type_cast_2664_wire;
      req <= phi_stmt_2658_req_0 & phi_stmt_2658_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2658",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2658_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2658,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2658
    phi_stmt_2665: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2668_wire & type_cast_2670_wire;
      req <= phi_stmt_2665_req_0 & phi_stmt_2665_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2665",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2665_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2665,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2665
    phi_stmt_2848: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2851_wire & type_cast_2854_wire_constant;
      req <= phi_stmt_2848_req_0 & phi_stmt_2848_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2848",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2848_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2848,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2848
    phi_stmt_2855: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2858_wire & type_cast_2860_wire;
      req <= phi_stmt_2855_req_0 & phi_stmt_2855_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2855",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2855_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2855,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2855
    phi_stmt_2861: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2864_wire & type_cast_2866_wire;
      req <= phi_stmt_2861_req_0 & phi_stmt_2861_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2861",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2861_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2861,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2861
    -- flow-through select operator MUX_2834_inst
    input_dim1x_x2_2835 <= type_cast_2832_wire_constant when (cmp111_2819(0) /=  '0') else inc_2814;
    addr_of_2750_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2750_final_reg_req_0;
      addr_of_2750_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2750_final_reg_req_1;
      addr_of_2750_final_reg_ack_1<= rack(0);
      addr_of_2750_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2750_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2749_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2773_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2773_final_reg_req_0;
      addr_of_2773_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2773_final_reg_req_1;
      addr_of_2773_final_reg_ack_1<= rack(0);
      addr_of_2773_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2773_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2772_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2774,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2561_inst_req_0;
      type_cast_2561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2561_inst_req_1;
      type_cast_2561_inst_ack_1<= rack(0);
      type_cast_2561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2574_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2574_inst_req_0;
      type_cast_2574_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2574_inst_req_1;
      type_cast_2574_inst_ack_1<= rack(0);
      type_cast_2574_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2574_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2571,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2575,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2632_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2632_inst_req_0;
      type_cast_2632_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2632_inst_req_1;
      type_cast_2632_inst_ack_1<= rack(0);
      type_cast_2632_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2632_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2589,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2633,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2636_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2636_inst_req_0;
      type_cast_2636_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2636_inst_req_1;
      type_cast_2636_inst_ack_1<= rack(0);
      type_cast_2636_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2636_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_2637,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2640_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2640_inst_req_0;
      type_cast_2640_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2640_inst_req_1;
      type_cast_2640_inst_ack_1<= rack(0);
      type_cast_2640_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2640_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_2641,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2650_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2650_inst_req_0;
      type_cast_2650_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2650_inst_req_1;
      type_cast_2650_inst_ack_1<= rack(0);
      type_cast_2650_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2650_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2873,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2650_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2657_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2657_inst_req_0;
      type_cast_2657_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2657_inst_req_1;
      type_cast_2657_inst_ack_1<= rack(0);
      type_cast_2657_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2657_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2848,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2657_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2664_inst_req_0;
      type_cast_2664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2664_inst_req_1;
      type_cast_2664_inst_ack_1<= rack(0);
      type_cast_2664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2855,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2664_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2668_inst_req_0;
      type_cast_2668_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2668_inst_req_1;
      type_cast_2668_inst_ack_1<= rack(0);
      type_cast_2668_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2668_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_2607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2668_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2670_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2670_inst_req_0;
      type_cast_2670_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2670_inst_req_1;
      type_cast_2670_inst_ack_1<= rack(0);
      type_cast_2670_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2670_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2861,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2670_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2705_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2705_inst_req_0;
      type_cast_2705_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2705_inst_req_1;
      type_cast_2705_inst_ack_1<= rack(0);
      type_cast_2705_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2705_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2651,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2709_inst_req_0;
      type_cast_2709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2709_inst_req_1;
      type_cast_2709_inst_ack_1<= rack(0);
      type_cast_2709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub67_2702,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2713_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2713_inst_req_0;
      type_cast_2713_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2713_inst_req_1;
      type_cast_2713_inst_ack_1<= rack(0);
      type_cast_2713_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2713_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub53_2692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2714,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2743_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2743_inst_req_0;
      type_cast_2743_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2743_inst_req_1;
      type_cast_2743_inst_ack_1<= rack(0);
      type_cast_2743_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2743_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr86_2740,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2744,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2781_inst_req_0;
      type_cast_2781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2781_inst_req_1;
      type_cast_2781_inst_ack_1<= rack(0);
      type_cast_2781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2781_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2651,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2822_inst_req_0;
      type_cast_2822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2822_inst_req_1;
      type_cast_2822_inst_ack_1<= rack(0);
      type_cast_2822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp111_2819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc115_2823,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2851_inst_req_0;
      type_cast_2851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2851_inst_req_1;
      type_cast_2851_inst_ack_1<= rack(0);
      type_cast_2851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add103_2806,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2851_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2858_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2858_inst_req_0;
      type_cast_2858_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2858_inst_req_1;
      type_cast_2858_inst_ack_1<= rack(0);
      type_cast_2858_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2858_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2658,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2858_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2860_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2860_inst_req_0;
      type_cast_2860_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2860_inst_req_1;
      type_cast_2860_inst_ack_1<= rack(0);
      type_cast_2860_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2860_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2835,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2860_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2864_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2864_inst_req_0;
      type_cast_2864_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2864_inst_req_1;
      type_cast_2864_inst_ack_1<= rack(0);
      type_cast_2864_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2864_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2864_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2866_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2866_inst_req_0;
      type_cast_2866_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2866_inst_req_1;
      type_cast_2866_inst_ack_1<= rack(0);
      type_cast_2866_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2866_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc115x_xinput_dim0x_x2_2828,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2866_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2749_index_1_rename
    process(R_idxprom_2748_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2748_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2748_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2749_index_1_resize
    process(idxprom_2744) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2744;
      ov := iv(13 downto 0);
      R_idxprom_2748_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2749_root_address_inst
    process(array_obj_ref_2749_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2749_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2749_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2772_index_1_rename
    process(R_idxprom91_2771_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom91_2771_resized;
      ov(13 downto 0) := iv;
      R_idxprom91_2771_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2772_index_1_resize
    process(idxprom91_2767) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom91_2767;
      ov := iv(13 downto 0);
      R_idxprom91_2771_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2772_root_address_inst
    process(array_obj_ref_2772_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2772_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2772_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2754_addr_0
    process(ptr_deref_2754_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2754_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2754_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2754_base_resize
    process(arrayidx87_2751) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2751;
      ov := iv(13 downto 0);
      ptr_deref_2754_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2754_gather_scatter
    process(ptr_deref_2754_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2754_data_0;
      ov(63 downto 0) := iv;
      tmp88_2755 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2754_root_address_inst
    process(ptr_deref_2754_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2754_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2754_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2776_addr_0
    process(ptr_deref_2776_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2776_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2776_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2776_base_resize
    process(arrayidx92_2774) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2774;
      ov := iv(13 downto 0);
      ptr_deref_2776_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2776_gather_scatter
    process(tmp88_2755) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp88_2755;
      ov(63 downto 0) := iv;
      ptr_deref_2776_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2776_root_address_inst
    process(ptr_deref_2776_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2776_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2776_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2794_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2793;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2794_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2794_branch_req_0,
          ack0 => if_stmt_2794_branch_ack_0,
          ack1 => if_stmt_2794_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2841_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp121_2840;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2841_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2841_branch_req_0,
          ack0 => if_stmt_2841_branch_ack_0,
          ack1 => if_stmt_2841_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2606_inst
    process(shr135_2596, shr31136_2602) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr135_2596, shr31136_2602, tmp_var);
      add32_2607 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2612_inst
    process(call7_2543) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2543, type_cast_2611_wire_constant, tmp_var);
      add50_2613 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2623_inst
    process(call9_2546) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2546, type_cast_2622_wire_constant, tmp_var);
      add63_2624 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2691_inst
    process(sub_2618, mul_2687) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2618, mul_2687, tmp_var);
      sub53_2692 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2701_inst
    process(sub66_2629, mul59_2697) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub66_2629, mul59_2697, tmp_var);
      sub67_2702 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2805_inst
    process(input_dim2x_x1_2651) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2651, type_cast_2804_wire_constant, tmp_var);
      add103_2806 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2813_inst
    process(input_dim1x_x1_2658) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2658, type_cast_2812_wire_constant, tmp_var);
      inc_2814 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2827_inst
    process(inc115_2823, input_dim0x_x2_2665) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc115_2823, input_dim0x_x2_2665, tmp_var);
      inc115x_xinput_dim0x_x2_2828 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2681_inst
    process(add_2580, tmp1_2677) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2580, tmp1_2677, tmp_var);
      add_src_0x_x0_2682 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2787_inst
    process(conv95_2782) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv95_2782, type_cast_2786_wire_constant, tmp_var);
      add96_2788 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2872_inst
    process(indvar_2644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2644, type_cast_2871_wire_constant, tmp_var);
      indvarx_xnext_2873 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2723_inst
    process(mul81_2719, conv75_2710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul81_2719, conv75_2710, tmp_var);
      add82_2724 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2733_inst
    process(mul83_2729, conv70_2706) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul83_2729, conv70_2706, tmp_var);
      add84_2734 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2766_inst
    process(shr90_2761) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr90_2761, type_cast_2765_wire_constant, tmp_var);
      idxprom91_2767 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2818_inst
    process(inc_2814, call1_2534) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2814, call1_2534, tmp_var);
      cmp111_2819 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2839_inst
    process(inc115x_xinput_dim0x_x2_2828, call_2531) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc115x_xinput_dim0x_x2_2828, call_2531, tmp_var);
      cmp121_2840 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2595_inst
    process(call_2531) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2531, type_cast_2594_wire_constant, tmp_var);
      shr135_2596 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2601_inst
    process(call_2531) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2531, type_cast_2600_wire_constant, tmp_var);
      shr31136_2602 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2739_inst
    process(add_src_0x_x0_2682) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2682, type_cast_2738_wire_constant, tmp_var);
      shr86_2740 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2760_inst
    process(add84_2734) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add84_2734, type_cast_2759_wire_constant, tmp_var);
      shr90_2761 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2686_inst
    process(input_dim0x_x2_2665, call13_2552) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2665, call13_2552, tmp_var);
      mul_2687 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2696_inst
    process(input_dim1x_x1_2658, call13_2552) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2658, call13_2552, tmp_var);
      mul59_2697 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2676_inst
    process(indvar_2644) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2644, type_cast_2675_wire_constant, tmp_var);
      tmp1_2677 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2718_inst
    process(conv80_2714, conv78_2637) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv80_2714, conv78_2637, tmp_var);
      mul81_2719 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2728_inst
    process(add82_2724, conv73_2633) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add82_2724, conv73_2633, tmp_var);
      mul83_2729 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2579_inst
    process(shl_2568, conv17_2575) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2568, conv17_2575, tmp_var);
      add_2580 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2567_inst
    process(conv_2562) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2562, type_cast_2566_wire_constant, tmp_var);
      shl_2568 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2617_inst
    process(add50_2613, call14_2555) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add50_2613, call14_2555, tmp_var);
      sub_2618 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2628_inst
    process(add63_2624, call14_2555) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add63_2624, call14_2555, tmp_var);
      sub66_2629 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2792_inst
    process(add96_2788, conv99_2641) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add96_2788, conv99_2641, tmp_var);
      cmp_2793 <= tmp_var; --
    end process;
    -- shared split operator group (30) : array_obj_ref_2749_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2748_scaled;
      array_obj_ref_2749_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2749_index_offset_req_0;
      array_obj_ref_2749_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2749_index_offset_req_1;
      array_obj_ref_2749_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_2772_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom91_2771_scaled;
      array_obj_ref_2772_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2772_index_offset_req_0;
      array_obj_ref_2772_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2772_index_offset_req_1;
      array_obj_ref_2772_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared load operator group (0) : ptr_deref_2754_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2754_load_0_req_0;
      ptr_deref_2754_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2754_load_0_req_1;
      ptr_deref_2754_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2754_word_address_0;
      ptr_deref_2754_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2776_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2776_store_0_req_0;
      ptr_deref_2776_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2776_store_0_req_1;
      ptr_deref_2776_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2776_word_address_0;
      data_in <= ptr_deref_2776_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2530_inst RPIPE_Block3_start_2533_inst RPIPE_Block3_start_2536_inst RPIPE_Block3_start_2539_inst RPIPE_Block3_start_2542_inst RPIPE_Block3_start_2545_inst RPIPE_Block3_start_2548_inst RPIPE_Block3_start_2551_inst RPIPE_Block3_start_2554_inst RPIPE_Block3_start_2557_inst RPIPE_Block3_start_2570_inst RPIPE_Block3_start_2582_inst RPIPE_Block3_start_2585_inst RPIPE_Block3_start_2588_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block3_start_2530_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_2533_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2536_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2539_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2542_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2545_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2548_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2551_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2554_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2557_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2570_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2582_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2585_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2588_inst_req_0;
      RPIPE_Block3_start_2530_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_2533_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2536_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2539_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2542_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2545_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2548_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2551_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2554_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2557_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2570_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2582_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2585_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2588_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block3_start_2530_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_2533_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2536_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2539_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2542_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2545_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2548_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2551_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2554_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2557_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2570_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2582_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2585_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2588_inst_req_1;
      RPIPE_Block3_start_2530_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_2533_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2536_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2539_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2542_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2545_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2548_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2551_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2554_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2557_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2570_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2582_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2585_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2588_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2531 <= data_out(223 downto 208);
      call1_2534 <= data_out(207 downto 192);
      call3_2537 <= data_out(191 downto 176);
      call5_2540 <= data_out(175 downto 160);
      call7_2543 <= data_out(159 downto 144);
      call9_2546 <= data_out(143 downto 128);
      call11_2549 <= data_out(127 downto 112);
      call13_2552 <= data_out(111 downto 96);
      call14_2555 <= data_out(95 downto 80);
      call15_2558 <= data_out(79 downto 64);
      call16_2571 <= data_out(63 downto 48);
      call18_2583 <= data_out(47 downto 32);
      call20_2586 <= data_out(31 downto 16);
      call22_2589 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2877_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2877_inst_req_0;
      WPIPE_Block3_done_2877_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2877_inst_req_1;
      WPIPE_Block3_done_2877_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2879_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_28_load_0_req_1 : boolean;
  signal LOAD_count_28_load_0_ack_1 : boolean;
  signal LOAD_count_28_load_0_req_0 : boolean;
  signal LOAD_count_28_load_0_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_29/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_sample_start_
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_update_start_
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/rr
      -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_28_load_0_req_1); -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_28_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_sample_completed_
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/ra
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_28_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/merge_ack
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_29/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_update_completed_
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_28_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_28_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_28_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_28_word_address_0 <= "0";
    -- equivalence LOAD_count_28_gather_scatter
    process(LOAD_count_28_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_28_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_28_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_28_load_0_req_0;
      LOAD_count_28_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_28_load_0_req_1;
      LOAD_count_28_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_28_word_address_0;
      LOAD_count_28_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(4 downto 4),
      memory_space_3_sr_ack => memory_space_3_sr_ack(4 downto 4),
      memory_space_3_sr_addr => memory_space_3_sr_addr(69 downto 56),
      memory_space_3_sr_data => memory_space_3_sr_data(319 downto 256),
      memory_space_3_sr_tag => memory_space_3_sr_tag(94 downto 76),
      memory_space_3_sc_req => memory_space_3_sc_req(4 downto 4),
      memory_space_3_sc_ack => memory_space_3_sc_ack(4 downto 4),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_sr_req => memory_space_3_sr_req(3 downto 3),
      memory_space_3_sr_ack => memory_space_3_sr_ack(3 downto 3),
      memory_space_3_sr_addr => memory_space_3_sr_addr(55 downto 42),
      memory_space_3_sr_data => memory_space_3_sr_data(255 downto 192),
      memory_space_3_sr_tag => memory_space_3_sr_tag(75 downto 57),
      memory_space_3_sc_req => memory_space_3_sc_req(3 downto 3),
      memory_space_3_sc_ack => memory_space_3_sc_ack(3 downto 3),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_sr_req => memory_space_3_sr_req(2 downto 2),
      memory_space_3_sr_ack => memory_space_3_sr_ack(2 downto 2),
      memory_space_3_sr_addr => memory_space_3_sr_addr(41 downto 28),
      memory_space_3_sr_data => memory_space_3_sr_data(191 downto 128),
      memory_space_3_sr_tag => memory_space_3_sr_tag(56 downto 38),
      memory_space_3_sc_req => memory_space_3_sc_req(2 downto 2),
      memory_space_3_sc_ack => memory_space_3_sc_ack(2 downto 2),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(37 downto 19),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
