-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    row_in : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
    input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_data : out  std_logic_vector(7 downto 0);
    input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_data : out  std_logic_vector(7 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(7 downto 0);
    input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe4_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 48)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal row_in_buffer :  std_logic_vector(15 downto 0);
  signal row_in_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal W_fetch_val2_322_delayed_13_0_340_inst_ack_0 : boolean;
  signal W_fetch_val2_322_delayed_13_0_340_inst_req_0 : boolean;
  signal W_fn2_320_delayed_13_0_337_inst_ack_1 : boolean;
  signal W_fetch_val2_322_delayed_13_0_340_inst_ack_1 : boolean;
  signal W_fetch_val2_322_delayed_13_0_340_inst_req_1 : boolean;
  signal W_fn2_320_delayed_13_0_337_inst_req_1 : boolean;
  signal W_fn2_314_delayed_7_0_329_inst_ack_0 : boolean;
  signal addr_of_327_final_reg_ack_1 : boolean;
  signal type_cast_371_inst_req_0 : boolean;
  signal addr_of_327_final_reg_req_1 : boolean;
  signal ptr_deref_335_load_0_ack_1 : boolean;
  signal ptr_deref_52_load_0_req_0 : boolean;
  signal ptr_deref_52_load_0_ack_0 : boolean;
  signal ptr_deref_263_load_0_ack_1 : boolean;
  signal ptr_deref_52_load_0_req_1 : boolean;
  signal ptr_deref_52_load_0_ack_1 : boolean;
  signal ptr_deref_335_load_0_req_1 : boolean;
  signal type_cast_299_inst_req_1 : boolean;
  signal array_obj_ref_75_index_offset_req_0 : boolean;
  signal array_obj_ref_75_index_offset_ack_0 : boolean;
  signal addr_of_327_final_reg_ack_0 : boolean;
  signal array_obj_ref_61_index_offset_req_0 : boolean;
  signal array_obj_ref_61_index_offset_ack_0 : boolean;
  signal W_fn2_320_delayed_13_0_337_inst_ack_0 : boolean;
  signal array_obj_ref_61_index_offset_req_1 : boolean;
  signal array_obj_ref_61_index_offset_ack_1 : boolean;
  signal W_fn2_314_delayed_7_0_329_inst_req_0 : boolean;
  signal addr_of_62_final_reg_req_0 : boolean;
  signal addr_of_62_final_reg_ack_0 : boolean;
  signal addr_of_62_final_reg_req_1 : boolean;
  signal addr_of_62_final_reg_ack_1 : boolean;
  signal ptr_deref_335_load_0_ack_0 : boolean;
  signal addr_of_327_final_reg_req_0 : boolean;
  signal W_fn2_320_delayed_13_0_337_inst_req_0 : boolean;
  signal ptr_deref_263_load_0_req_1 : boolean;
  signal ptr_deref_66_load_0_req_0 : boolean;
  signal ptr_deref_66_load_0_ack_0 : boolean;
  signal ptr_deref_66_load_0_req_1 : boolean;
  signal ptr_deref_66_load_0_ack_1 : boolean;
  signal ptr_deref_335_load_0_req_0 : boolean;
  signal type_cast_299_inst_ack_1 : boolean;
  signal phi_stmt_102_ack_0 : boolean;
  signal array_obj_ref_75_index_offset_req_1 : boolean;
  signal array_obj_ref_75_index_offset_ack_1 : boolean;
  signal addr_of_76_final_reg_req_0 : boolean;
  signal addr_of_76_final_reg_ack_0 : boolean;
  signal addr_of_76_final_reg_req_1 : boolean;
  signal addr_of_76_final_reg_ack_1 : boolean;
  signal addr_of_255_final_reg_ack_0 : boolean;
  signal ptr_deref_80_load_0_req_0 : boolean;
  signal type_cast_299_inst_ack_0 : boolean;
  signal ptr_deref_80_load_0_ack_0 : boolean;
  signal addr_of_255_final_reg_ack_1 : boolean;
  signal ptr_deref_263_load_0_ack_0 : boolean;
  signal ptr_deref_80_load_0_req_1 : boolean;
  signal ptr_deref_80_load_0_ack_1 : boolean;
  signal type_cast_299_inst_req_0 : boolean;
  signal array_obj_ref_93_index_offset_req_0 : boolean;
  signal array_obj_ref_93_index_offset_ack_0 : boolean;
  signal array_obj_ref_93_index_offset_req_1 : boolean;
  signal array_obj_ref_93_index_offset_ack_1 : boolean;
  signal addr_of_94_final_reg_req_0 : boolean;
  signal addr_of_94_final_reg_ack_0 : boolean;
  signal addr_of_94_final_reg_req_1 : boolean;
  signal addr_of_94_final_reg_ack_1 : boolean;
  signal array_obj_ref_326_index_offset_ack_1 : boolean;
  signal array_obj_ref_326_index_offset_req_1 : boolean;
  signal ptr_deref_263_load_0_req_0 : boolean;
  signal ptr_deref_98_load_0_req_0 : boolean;
  signal ptr_deref_98_load_0_ack_0 : boolean;
  signal addr_of_255_final_reg_req_1 : boolean;
  signal ptr_deref_98_load_0_req_1 : boolean;
  signal ptr_deref_98_load_0_ack_1 : boolean;
  signal do_while_stmt_100_branch_req_0 : boolean;
  signal addr_of_255_final_reg_req_0 : boolean;
  signal phi_stmt_102_req_1 : boolean;
  signal phi_stmt_102_req_0 : boolean;
  signal n_fetch_val1_276_132_buf_req_0 : boolean;
  signal n_fetch_val1_276_132_buf_ack_0 : boolean;
  signal n_fetch_val1_276_132_buf_req_1 : boolean;
  signal n_fetch_val1_276_132_buf_ack_1 : boolean;
  signal n_address1_236_106_buf_req_0 : boolean;
  signal n_address1_236_106_buf_ack_0 : boolean;
  signal n_address1_236_106_buf_req_1 : boolean;
  signal n_address1_236_106_buf_ack_1 : boolean;
  signal phi_stmt_107_req_1 : boolean;
  signal phi_stmt_107_req_0 : boolean;
  signal phi_stmt_107_ack_0 : boolean;
  signal type_cast_110_inst_req_0 : boolean;
  signal type_cast_110_inst_ack_0 : boolean;
  signal type_cast_110_inst_req_1 : boolean;
  signal type_cast_110_inst_ack_1 : boolean;
  signal array_obj_ref_326_index_offset_ack_0 : boolean;
  signal W_fetch_val1_262_delayed_13_0_268_inst_ack_1 : boolean;
  signal W_fetch_val1_262_delayed_13_0_268_inst_req_1 : boolean;
  signal n_address2_308_111_buf_req_0 : boolean;
  signal n_address2_308_111_buf_ack_0 : boolean;
  signal n_address2_308_111_buf_req_1 : boolean;
  signal n_address2_308_111_buf_ack_1 : boolean;
  signal W_fetch_val1_262_delayed_13_0_268_inst_ack_0 : boolean;
  signal W_fetch_val1_262_delayed_13_0_268_inst_req_0 : boolean;
  signal phi_stmt_112_req_1 : boolean;
  signal phi_stmt_112_req_0 : boolean;
  signal phi_stmt_112_ack_0 : boolean;
  signal type_cast_115_inst_req_0 : boolean;
  signal type_cast_115_inst_ack_0 : boolean;
  signal type_cast_115_inst_req_1 : boolean;
  signal type_cast_115_inst_ack_1 : boolean;
  signal n_address3_380_116_buf_req_0 : boolean;
  signal n_address3_380_116_buf_ack_0 : boolean;
  signal W_fn1_254_delayed_7_0_257_inst_ack_1 : boolean;
  signal W_fn1_254_delayed_7_0_257_inst_req_1 : boolean;
  signal n_address3_380_116_buf_req_1 : boolean;
  signal n_address3_380_116_buf_ack_1 : boolean;
  signal phi_stmt_117_req_1 : boolean;
  signal phi_stmt_117_req_0 : boolean;
  signal phi_stmt_117_ack_0 : boolean;
  signal W_fn1_260_delayed_13_0_265_inst_ack_1 : boolean;
  signal W_fn1_260_delayed_13_0_265_inst_req_1 : boolean;
  signal W_fn2_314_delayed_7_0_329_inst_ack_1 : boolean;
  signal type_cast_122_inst_req_0 : boolean;
  signal type_cast_122_inst_ack_0 : boolean;
  signal type_cast_122_inst_req_1 : boolean;
  signal type_cast_122_inst_ack_1 : boolean;
  signal W_fn1_254_delayed_7_0_257_inst_ack_0 : boolean;
  signal array_obj_ref_326_index_offset_req_0 : boolean;
  signal W_fn1_254_delayed_7_0_257_inst_req_0 : boolean;
  signal W_fn1_260_delayed_13_0_265_inst_ack_0 : boolean;
  signal W_fn1_260_delayed_13_0_265_inst_req_0 : boolean;
  signal W_fn2_314_delayed_7_0_329_inst_req_1 : boolean;
  signal n_address4_452_123_buf_req_0 : boolean;
  signal n_address4_452_123_buf_ack_0 : boolean;
  signal n_address4_452_123_buf_req_1 : boolean;
  signal n_address4_452_123_buf_ack_1 : boolean;
  signal phi_stmt_124_req_1 : boolean;
  signal phi_stmt_124_req_0 : boolean;
  signal phi_stmt_124_ack_0 : boolean;
  signal n_mycounter_168_128_buf_req_0 : boolean;
  signal n_mycounter_168_128_buf_ack_0 : boolean;
  signal n_mycounter_168_128_buf_req_1 : boolean;
  signal n_mycounter_168_128_buf_ack_1 : boolean;
  signal phi_stmt_129_req_1 : boolean;
  signal phi_stmt_129_req_0 : boolean;
  signal phi_stmt_129_ack_0 : boolean;
  signal my_fetch1_53_131_buf_req_0 : boolean;
  signal my_fetch1_53_131_buf_ack_0 : boolean;
  signal my_fetch1_53_131_buf_req_1 : boolean;
  signal my_fetch1_53_131_buf_ack_1 : boolean;
  signal phi_stmt_133_req_1 : boolean;
  signal phi_stmt_133_req_0 : boolean;
  signal phi_stmt_133_ack_0 : boolean;
  signal my_fetch2_67_135_buf_req_0 : boolean;
  signal my_fetch2_67_135_buf_ack_0 : boolean;
  signal my_fetch2_67_135_buf_req_1 : boolean;
  signal my_fetch2_67_135_buf_ack_1 : boolean;
  signal type_cast_371_inst_ack_0 : boolean;
  signal type_cast_371_inst_req_1 : boolean;
  signal n_fetch_val2_348_136_buf_req_0 : boolean;
  signal n_fetch_val2_348_136_buf_ack_0 : boolean;
  signal n_fetch_val2_348_136_buf_req_1 : boolean;
  signal n_fetch_val2_348_136_buf_ack_1 : boolean;
  signal phi_stmt_137_req_1 : boolean;
  signal phi_stmt_137_req_0 : boolean;
  signal phi_stmt_137_ack_0 : boolean;
  signal my_fetch3_81_139_buf_req_0 : boolean;
  signal my_fetch3_81_139_buf_ack_0 : boolean;
  signal my_fetch3_81_139_buf_req_1 : boolean;
  signal my_fetch3_81_139_buf_ack_1 : boolean;
  signal n_fetch_val3_420_140_buf_req_0 : boolean;
  signal n_fetch_val3_420_140_buf_ack_0 : boolean;
  signal n_fetch_val3_420_140_buf_req_1 : boolean;
  signal n_fetch_val3_420_140_buf_ack_1 : boolean;
  signal phi_stmt_141_req_1 : boolean;
  signal phi_stmt_141_req_0 : boolean;
  signal phi_stmt_141_ack_0 : boolean;
  signal my_fetch4_99_143_buf_req_0 : boolean;
  signal my_fetch4_99_143_buf_ack_0 : boolean;
  signal my_fetch4_99_143_buf_req_1 : boolean;
  signal my_fetch4_99_143_buf_ack_1 : boolean;
  signal n_fetch_val4_492_144_buf_req_0 : boolean;
  signal n_fetch_val4_492_144_buf_ack_0 : boolean;
  signal n_fetch_val4_492_144_buf_req_1 : boolean;
  signal n_fetch_val4_492_144_buf_ack_1 : boolean;
  signal phi_stmt_145_req_1 : boolean;
  signal phi_stmt_145_req_0 : boolean;
  signal phi_stmt_145_ack_0 : boolean;
  signal n_row1_186_149_buf_req_0 : boolean;
  signal n_row1_186_149_buf_ack_0 : boolean;
  signal n_row1_186_149_buf_req_1 : boolean;
  signal n_row1_186_149_buf_ack_1 : boolean;
  signal phi_stmt_150_req_1 : boolean;
  signal phi_stmt_150_req_0 : boolean;
  signal phi_stmt_150_ack_0 : boolean;
  signal n_row2_194_154_buf_req_0 : boolean;
  signal n_row2_194_154_buf_ack_0 : boolean;
  signal n_row2_194_154_buf_req_1 : boolean;
  signal n_row2_194_154_buf_ack_1 : boolean;
  signal type_cast_227_inst_req_0 : boolean;
  signal type_cast_227_inst_ack_0 : boolean;
  signal type_cast_227_inst_req_1 : boolean;
  signal type_cast_227_inst_ack_1 : boolean;
  signal array_obj_ref_254_index_offset_req_0 : boolean;
  signal array_obj_ref_254_index_offset_ack_0 : boolean;
  signal array_obj_ref_254_index_offset_req_1 : boolean;
  signal array_obj_ref_254_index_offset_ack_1 : boolean;
  signal type_cast_371_inst_ack_1 : boolean;
  signal array_obj_ref_398_index_offset_req_0 : boolean;
  signal array_obj_ref_398_index_offset_ack_0 : boolean;
  signal array_obj_ref_398_index_offset_req_1 : boolean;
  signal array_obj_ref_398_index_offset_ack_1 : boolean;
  signal addr_of_399_final_reg_req_0 : boolean;
  signal addr_of_399_final_reg_ack_0 : boolean;
  signal addr_of_399_final_reg_req_1 : boolean;
  signal addr_of_399_final_reg_ack_1 : boolean;
  signal W_fn3_374_delayed_7_0_401_inst_req_0 : boolean;
  signal W_fn3_374_delayed_7_0_401_inst_ack_0 : boolean;
  signal W_fn3_374_delayed_7_0_401_inst_req_1 : boolean;
  signal W_fn3_374_delayed_7_0_401_inst_ack_1 : boolean;
  signal ptr_deref_407_load_0_req_0 : boolean;
  signal ptr_deref_407_load_0_ack_0 : boolean;
  signal ptr_deref_407_load_0_req_1 : boolean;
  signal ptr_deref_407_load_0_ack_1 : boolean;
  signal W_fn3_380_delayed_13_0_409_inst_req_0 : boolean;
  signal W_fn3_380_delayed_13_0_409_inst_ack_0 : boolean;
  signal W_fn3_380_delayed_13_0_409_inst_req_1 : boolean;
  signal W_fn3_380_delayed_13_0_409_inst_ack_1 : boolean;
  signal W_fetch_val3_382_delayed_13_0_412_inst_req_0 : boolean;
  signal W_fetch_val3_382_delayed_13_0_412_inst_ack_0 : boolean;
  signal W_fetch_val3_382_delayed_13_0_412_inst_req_1 : boolean;
  signal W_fetch_val3_382_delayed_13_0_412_inst_ack_1 : boolean;
  signal type_cast_443_inst_req_0 : boolean;
  signal type_cast_443_inst_ack_0 : boolean;
  signal type_cast_443_inst_req_1 : boolean;
  signal type_cast_443_inst_ack_1 : boolean;
  signal array_obj_ref_470_index_offset_req_0 : boolean;
  signal array_obj_ref_470_index_offset_ack_0 : boolean;
  signal array_obj_ref_470_index_offset_req_1 : boolean;
  signal array_obj_ref_470_index_offset_ack_1 : boolean;
  signal addr_of_471_final_reg_req_0 : boolean;
  signal addr_of_471_final_reg_ack_0 : boolean;
  signal addr_of_471_final_reg_req_1 : boolean;
  signal addr_of_471_final_reg_ack_1 : boolean;
  signal W_fn4_434_delayed_7_0_473_inst_req_0 : boolean;
  signal W_fn4_434_delayed_7_0_473_inst_ack_0 : boolean;
  signal W_fn4_434_delayed_7_0_473_inst_req_1 : boolean;
  signal W_fn4_434_delayed_7_0_473_inst_ack_1 : boolean;
  signal ptr_deref_479_load_0_req_0 : boolean;
  signal ptr_deref_479_load_0_ack_0 : boolean;
  signal ptr_deref_479_load_0_req_1 : boolean;
  signal ptr_deref_479_load_0_ack_1 : boolean;
  signal W_fn4_440_delayed_13_0_481_inst_req_0 : boolean;
  signal W_fn4_440_delayed_13_0_481_inst_ack_0 : boolean;
  signal W_fn4_440_delayed_13_0_481_inst_req_1 : boolean;
  signal W_fn4_440_delayed_13_0_481_inst_ack_1 : boolean;
  signal W_fetch_val4_442_delayed_13_0_484_inst_req_0 : boolean;
  signal W_fetch_val4_442_delayed_13_0_484_inst_ack_0 : boolean;
  signal W_fetch_val4_442_delayed_13_0_484_inst_req_1 : boolean;
  signal W_fetch_val4_442_delayed_13_0_484_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_494_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_494_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_494_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_494_inst_ack_1 : boolean;
  signal WPIPE_input_pipe2_498_inst_req_0 : boolean;
  signal WPIPE_input_pipe2_498_inst_ack_0 : boolean;
  signal WPIPE_input_pipe2_498_inst_req_1 : boolean;
  signal WPIPE_input_pipe2_498_inst_ack_1 : boolean;
  signal WPIPE_input_pipe3_502_inst_req_0 : boolean;
  signal WPIPE_input_pipe3_502_inst_ack_0 : boolean;
  signal WPIPE_input_pipe3_502_inst_req_1 : boolean;
  signal WPIPE_input_pipe3_502_inst_ack_1 : boolean;
  signal WPIPE_input_pipe4_506_inst_req_0 : boolean;
  signal WPIPE_input_pipe4_506_inst_ack_0 : boolean;
  signal WPIPE_input_pipe4_506_inst_req_1 : boolean;
  signal WPIPE_input_pipe4_506_inst_ack_1 : boolean;
  signal do_while_stmt_100_branch_ack_0 : boolean;
  signal do_while_stmt_100_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 48) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= row_in;
  row_in_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= ct;
  ct_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(tag_length + 47 downto 48) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 47 downto 48);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(377 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0:  members (103) 
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_29/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/branch_block_stmt_29__entry__
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99__entry__
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_update_start
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_resized_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_scaled_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_computed_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_resize_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_resize_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_resize_1/index_resize_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_scale_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_scale_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_update_start
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_complete/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_resized_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_scaled_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_computed_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_resize_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_resize_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_resize_1/index_resize_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_scale_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_scale_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_complete/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_resized_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_scaled_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_computed_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_resize_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_resize_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_resize_1/index_resize_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_scale_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_scale_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_update_start
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_complete/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/word_0/cr
      -- 
    rr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_52_load_0_req_0); -- 
    cr_58_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_58_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_52_load_0_req_1); -- 
    req_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_75_index_offset_req_0); -- 
    req_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_61_index_offset_req_0); -- 
    req_94_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_94_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_61_index_offset_req_1); -- 
    req_109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => addr_of_62_final_reg_req_1); -- 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_66_load_0_req_1); -- 
    req_190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_75_index_offset_req_1); -- 
    req_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => addr_of_76_final_reg_req_1); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_80_load_0_req_1); -- 
    req_281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_93_index_offset_req_0); -- 
    req_286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_93_index_offset_req_1); -- 
    req_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => addr_of_94_final_reg_req_1); -- 
    cr_346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_98_load_0_req_1); -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	377 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_29/do_while_stmt_100__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_29/$exit
      -- CP-element group 1: 	 branch_block_stmt_29/branch_block_stmt_29__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(377);
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/$exit
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/word_0/ra
      -- 
    ra_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_52_load_0_ack_0, ack => access_T_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	22 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/$exit
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/word_0/ca
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/ptr_deref_52_Merge/$entry
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/ptr_deref_52_Merge/$exit
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/ptr_deref_52_Merge/merge_req
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/ptr_deref_52_Merge/merge_ack
      -- 
    ca_59_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_52_load_0_ack_1, ack => access_T_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	22 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_sample_complete
      -- CP-element group 4: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Sample/ack
      -- 
    ack_90_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_61_index_offset_ack_0, ack => access_T_CP_0_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (11) 
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_root_address_calculated
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_offset_calculated
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Update/ack
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_base_plus_offset/$entry
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_base_plus_offset/$exit
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_base_plus_offset/sum_rename_req
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_base_plus_offset/sum_rename_ack
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_request/$entry
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_request/req
      -- 
    ack_95_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_61_index_offset_ack_1, ack => access_T_CP_0_elements(5)); -- 
    req_104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(5), ack => addr_of_62_final_reg_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_request/$exit
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_request/ack
      -- 
    ack_105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_62_final_reg_ack_0, ack => access_T_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (24) 
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_complete/ack
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_word_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_root_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_address_resized
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_addr_resize/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_addr_resize/$exit
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_addr_resize/base_resize_req
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_addr_resize/base_resize_ack
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_plus_offset/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_plus_offset/$exit
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_plus_offset/sum_rename_req
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_plus_offset/sum_rename_ack
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_word_addrgen/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_word_addrgen/$exit
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_word_addrgen/root_register_req
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_word_addrgen/root_register_ack
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/word_0/rr
      -- 
    ack_110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_62_final_reg_ack_1, ack => access_T_CP_0_elements(7)); -- 
    rr_143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(7), ack => ptr_deref_66_load_0_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/$exit
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/word_0/ra
      -- 
    ra_144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_66_load_0_ack_0, ack => access_T_CP_0_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	22 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/ptr_deref_66_Merge/$entry
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/ptr_deref_66_Merge/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/ptr_deref_66_Merge/merge_req
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/ptr_deref_66_Merge/merge_ack
      -- 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_66_load_0_ack_1, ack => access_T_CP_0_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	22 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_sample_complete
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Sample/ack
      -- 
    ack_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_75_index_offset_ack_0, ack => access_T_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (11) 
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_offset_calculated
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Update/ack
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_base_plus_offset/$entry
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_base_plus_offset/$exit
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_base_plus_offset/sum_rename_req
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_base_plus_offset/sum_rename_ack
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_request/$entry
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_request/req
      -- 
    ack_191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_75_index_offset_ack_1, ack => access_T_CP_0_elements(11)); -- 
    req_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(11), ack => addr_of_76_final_reg_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_request/$exit
      -- CP-element group 12: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_request/ack
      -- 
    ack_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_76_final_reg_ack_0, ack => access_T_CP_0_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (24) 
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_complete/ack
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_word_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_address_resized
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_addr_resize/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_addr_resize/$exit
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_addr_resize/base_resize_req
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_addr_resize/base_resize_ack
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_word_addrgen/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_word_addrgen/$exit
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_word_addrgen/root_register_req
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_word_addrgen/root_register_ack
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/word_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/word_0/rr
      -- 
    ack_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_76_final_reg_ack_1, ack => access_T_CP_0_elements(13)); -- 
    rr_239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(13), ack => ptr_deref_80_load_0_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/$exit
      -- CP-element group 14: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/word_0/ra
      -- 
    ra_240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_80_load_0_ack_0, ack => access_T_CP_0_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	22 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/word_0/ca
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/ptr_deref_80_Merge/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/ptr_deref_80_Merge/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/ptr_deref_80_Merge/merge_req
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/ptr_deref_80_Merge/merge_ack
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_80_load_0_ack_1, ack => access_T_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_sample_complete
      -- CP-element group 16: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Sample/ack
      -- 
    ack_282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_93_index_offset_ack_0, ack => access_T_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (11) 
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_root_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_offset_calculated
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Update/ack
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_base_plus_offset/$entry
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_base_plus_offset/$exit
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_base_plus_offset/sum_rename_req
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_base_plus_offset/sum_rename_ack
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_request/$entry
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_request/req
      -- 
    ack_287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_93_index_offset_ack_1, ack => access_T_CP_0_elements(17)); -- 
    req_296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(17), ack => addr_of_94_final_reg_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_request/$exit
      -- CP-element group 18: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_request/ack
      -- 
    ack_297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_94_final_reg_ack_0, ack => access_T_CP_0_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (24) 
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_complete/$exit
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_complete/ack
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_word_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_root_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_address_resized
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_addr_resize/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_addr_resize/$exit
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_addr_resize/base_resize_req
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_addr_resize/base_resize_ack
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_plus_offset/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_plus_offset/$exit
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_plus_offset/sum_rename_ack
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_word_addrgen/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_word_addrgen/$exit
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_word_addrgen/root_register_req
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_word_addrgen/root_register_ack
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/word_0/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/word_0/rr
      -- 
    ack_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_94_final_reg_ack_1, ack => access_T_CP_0_elements(19)); -- 
    rr_335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(19), ack => ptr_deref_98_load_0_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/word_0/ra
      -- 
    ra_336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_98_load_0_ack_0, ack => access_T_CP_0_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/word_0/ca
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/ptr_deref_98_Merge/$entry
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/ptr_deref_98_Merge/$exit
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/ptr_deref_98_Merge/merge_req
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/ptr_deref_98_Merge/merge_ack
      -- 
    ca_347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_98_load_0_ack_1, ack => access_T_CP_0_elements(21)); -- 
    -- CP-element group 22:  join  transition  place  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: 	16 
    -- CP-element group 22: 	3 
    -- CP-element group 22: 	4 
    -- CP-element group 22: 	9 
    -- CP-element group 22: 	10 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99__exit__
      -- CP-element group 22: 	 branch_block_stmt_29/do_while_stmt_100__entry__
      -- CP-element group 22: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/$exit
      -- 
    access_T_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(21) & access_T_CP_0_elements(16) & access_T_CP_0_elements(3) & access_T_CP_0_elements(4) & access_T_CP_0_elements(9) & access_T_CP_0_elements(10) & access_T_CP_0_elements(15);
      gj_access_T_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  place  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	29 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_29/do_while_stmt_100/$entry
      -- CP-element group 23: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100__entry__
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(22);
    -- CP-element group 24:  merge  place  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	377 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100__exit__
      -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  merge  place  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_29/do_while_stmt_100/loop_back
      -- 
    -- Element group access_T_CP_0_elements(25) is bound as output of CP function.
    -- CP-element group 26:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	375 
    -- CP-element group 26: 	376 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_100/condition_done
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_100/loop_exit/$entry
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_100/loop_taken/$entry
      -- 
    access_T_CP_0_elements(26) <= access_T_CP_0_elements(31);
    -- CP-element group 27:  branch  place  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	374 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_29/do_while_stmt_100/loop_body_done
      -- 
    access_T_CP_0_elements(27) <= access_T_CP_0_elements(374);
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	141 
    -- CP-element group 28: 	160 
    -- CP-element group 28: 	42 
    -- CP-element group 28: 	82 
    -- CP-element group 28: 	124 
    -- CP-element group 28: 	103 
    -- CP-element group 28: 	61 
    -- CP-element group 28: 	179 
    -- CP-element group 28: 	198 
    -- CP-element group 28: 	217 
    -- CP-element group 28: 	236 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(28) <= access_T_CP_0_elements(25);
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	143 
    -- CP-element group 29: 	162 
    -- CP-element group 29: 	84 
    -- CP-element group 29: 	126 
    -- CP-element group 29: 	44 
    -- CP-element group 29: 	105 
    -- CP-element group 29: 	63 
    -- CP-element group 29: 	181 
    -- CP-element group 29: 	200 
    -- CP-element group 29: 	219 
    -- CP-element group 29: 	238 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(29) <= access_T_CP_0_elements(23);
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	137 
    -- CP-element group 30: 	138 
    -- CP-element group 30: 	154 
    -- CP-element group 30: 	155 
    -- CP-element group 30: 	173 
    -- CP-element group 30: 	36 
    -- CP-element group 30: 	55 
    -- CP-element group 30: 	56 
    -- CP-element group 30: 	76 
    -- CP-element group 30: 	77 
    -- CP-element group 30: 	37 
    -- CP-element group 30: 	118 
    -- CP-element group 30: 	119 
    -- CP-element group 30: 	97 
    -- CP-element group 30: 	98 
    -- CP-element group 30: 	174 
    -- CP-element group 30: 	192 
    -- CP-element group 30: 	193 
    -- CP-element group 30: 	211 
    -- CP-element group 30: 	212 
    -- CP-element group 30: 	230 
    -- CP-element group 30: 	231 
    -- CP-element group 30: 	249 
    -- CP-element group 30: 	254 
    -- CP-element group 30: 	256 
    -- CP-element group 30: 	277 
    -- CP-element group 30: 	282 
    -- CP-element group 30: 	284 
    -- CP-element group 30: 	305 
    -- CP-element group 30: 	310 
    -- CP-element group 30: 	312 
    -- CP-element group 30: 	333 
    -- CP-element group 30: 	338 
    -- CP-element group 30: 	340 
    -- CP-element group 30: 	373 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/$entry
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	35 
    -- CP-element group 31: 	123 
    -- CP-element group 31: 	216 
    -- CP-element group 31: 	373 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	26 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/condition_evaluated
      -- 
    condition_evaluated_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(31), ack => do_while_stmt_100_branch_req_0); -- 
    access_T_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(35) & access_T_CP_0_elements(123) & access_T_CP_0_elements(216) & access_T_CP_0_elements(373);
      gj_access_T_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	137 
    -- CP-element group 32: 	154 
    -- CP-element group 32: 	173 
    -- CP-element group 32: 	36 
    -- CP-element group 32: 	55 
    -- CP-element group 32: 	76 
    -- CP-element group 32: 	118 
    -- CP-element group 32: 	97 
    -- CP-element group 32: 	192 
    -- CP-element group 32: 	211 
    -- CP-element group 32: 	230 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	35 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	156 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	78 
    -- CP-element group 32: 	120 
    -- CP-element group 32: 	99 
    -- CP-element group 32: 	38 
    -- CP-element group 32: 	175 
    -- CP-element group 32: 	194 
    -- CP-element group 32: 	213 
    -- CP-element group 32: 	232 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/aggregated_phi_sample_req
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_sample_start__ps
      -- 
    access_T_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= access_T_CP_0_elements(137) & access_T_CP_0_elements(154) & access_T_CP_0_elements(173) & access_T_CP_0_elements(36) & access_T_CP_0_elements(55) & access_T_CP_0_elements(76) & access_T_CP_0_elements(118) & access_T_CP_0_elements(97) & access_T_CP_0_elements(192) & access_T_CP_0_elements(211) & access_T_CP_0_elements(230) & access_T_CP_0_elements(35);
      gj_access_T_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	139 
    -- CP-element group 33: 	157 
    -- CP-element group 33: 	58 
    -- CP-element group 33: 	79 
    -- CP-element group 33: 	121 
    -- CP-element group 33: 	100 
    -- CP-element group 33: 	39 
    -- CP-element group 33: 	176 
    -- CP-element group 33: 	195 
    -- CP-element group 33: 	214 
    -- CP-element group 33: 	233 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	250 
    -- CP-element group 33: 	266 
    -- CP-element group 33: 	270 
    -- CP-element group 33: 	274 
    -- CP-element group 33: 	278 
    -- CP-element group 33: 	294 
    -- CP-element group 33: 	298 
    -- CP-element group 33: 	302 
    -- CP-element group 33: 	306 
    -- CP-element group 33: 	322 
    -- CP-element group 33: 	326 
    -- CP-element group 33: 	330 
    -- CP-element group 33: 	334 
    -- CP-element group 33: 	350 
    -- CP-element group 33: 	354 
    -- CP-element group 33: 	358 
    -- CP-element group 33: 	374 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	137 
    -- CP-element group 33: 	154 
    -- CP-element group 33: 	173 
    -- CP-element group 33: 	36 
    -- CP-element group 33: 	55 
    -- CP-element group 33: 	76 
    -- CP-element group 33: 	118 
    -- CP-element group 33: 	97 
    -- CP-element group 33: 	192 
    -- CP-element group 33: 	211 
    -- CP-element group 33: 	230 
    -- CP-element group 33:  members (12) 
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/aggregated_phi_sample_ack
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_sample_completed_
      -- 
    access_T_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= access_T_CP_0_elements(139) & access_T_CP_0_elements(157) & access_T_CP_0_elements(58) & access_T_CP_0_elements(79) & access_T_CP_0_elements(121) & access_T_CP_0_elements(100) & access_T_CP_0_elements(39) & access_T_CP_0_elements(176) & access_T_CP_0_elements(195) & access_T_CP_0_elements(214) & access_T_CP_0_elements(233);
      gj_access_T_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	138 
    -- CP-element group 34: 	155 
    -- CP-element group 34: 	56 
    -- CP-element group 34: 	77 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	119 
    -- CP-element group 34: 	98 
    -- CP-element group 34: 	174 
    -- CP-element group 34: 	193 
    -- CP-element group 34: 	212 
    -- CP-element group 34: 	231 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	158 
    -- CP-element group 34: 	59 
    -- CP-element group 34: 	80 
    -- CP-element group 34: 	122 
    -- CP-element group 34: 	101 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	177 
    -- CP-element group 34: 	196 
    -- CP-element group 34: 	215 
    -- CP-element group 34: 	234 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/aggregated_phi_update_req
      -- CP-element group 34: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_update_start__ps
      -- 
    access_T_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= access_T_CP_0_elements(138) & access_T_CP_0_elements(155) & access_T_CP_0_elements(56) & access_T_CP_0_elements(77) & access_T_CP_0_elements(37) & access_T_CP_0_elements(119) & access_T_CP_0_elements(98) & access_T_CP_0_elements(174) & access_T_CP_0_elements(193) & access_T_CP_0_elements(212) & access_T_CP_0_elements(231);
      gj_access_T_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	140 
    -- CP-element group 35: 	159 
    -- CP-element group 35: 	60 
    -- CP-element group 35: 	41 
    -- CP-element group 35: 	81 
    -- CP-element group 35: 	123 
    -- CP-element group 35: 	102 
    -- CP-element group 35: 	178 
    -- CP-element group 35: 	197 
    -- CP-element group 35: 	216 
    -- CP-element group 35: 	235 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	31 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	32 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= access_T_CP_0_elements(140) & access_T_CP_0_elements(159) & access_T_CP_0_elements(60) & access_T_CP_0_elements(41) & access_T_CP_0_elements(81) & access_T_CP_0_elements(123) & access_T_CP_0_elements(102) & access_T_CP_0_elements(178) & access_T_CP_0_elements(197) & access_T_CP_0_elements(216) & access_T_CP_0_elements(235);
      gj_access_T_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	30 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: 	252 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	32 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_sample_start_
      -- 
    access_T_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(252);
      gj_access_T_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	30 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	41 
    -- CP-element group 37: 	257 
    -- CP-element group 37: 	263 
    -- CP-element group 37: 	271 
    -- CP-element group 37: 	362 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	34 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_update_start_
      -- 
    access_T_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(41) & access_T_CP_0_elements(257) & access_T_CP_0_elements(263) & access_T_CP_0_elements(271) & access_T_CP_0_elements(362);
      gj_access_T_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	32 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_sample_start__ps
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(32);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	33 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_update_start__ps
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(34);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	35 
    -- CP-element group 41: 	255 
    -- CP-element group 41: 	261 
    -- CP-element group 41: 	269 
    -- CP-element group 41: 	361 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	37 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	28 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_loopback_trigger
      -- 
    access_T_CP_0_elements(42) <= access_T_CP_0_elements(28);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_loopback_sample_req
      -- CP-element group 43: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_loopback_sample_req_ps
      -- 
    phi_stmt_102_loopback_sample_req_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_102_loopback_sample_req_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => phi_stmt_102_req_1); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	29 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_entry_trigger
      -- 
    access_T_CP_0_elements(44) <= access_T_CP_0_elements(29);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_entry_sample_req
      -- CP-element group 45: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_entry_sample_req_ps
      -- 
    phi_stmt_102_entry_sample_req_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_102_entry_sample_req_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(45), ack => phi_stmt_102_req_0); -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_phi_mux_ack
      -- CP-element group 46: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_phi_mux_ack_ps
      -- 
    phi_stmt_102_phi_mux_ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_102_ack_0, ack => access_T_CP_0_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_sample_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_update_start_
      -- 
    -- Element group access_T_CP_0_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_update_completed__ps
      -- 
    access_T_CP_0_elements(49) <= access_T_CP_0_elements(50);
    -- CP-element group 50:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	49 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(48), ack => access_T_CP_0_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_sample_start__ps
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Sample/req
      -- 
    req_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(51), ack => n_address1_236_106_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_update_start__ps
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_update_start_
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Update/req
      -- 
    req_414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(52), ack => n_address1_236_106_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Sample/ack
      -- 
    ack_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_236_106_buf_ack_0, ack => access_T_CP_0_elements(53)); -- 
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Update/ack
      -- 
    ack_415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_236_106_buf_ack_1, ack => access_T_CP_0_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	30 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	33 
    -- CP-element group 55: 	280 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	32 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_sample_start_
      -- 
    access_T_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(280);
      gj_access_T_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	30 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	285 
    -- CP-element group 56: 	291 
    -- CP-element group 56: 	299 
    -- CP-element group 56: 	365 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	34 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_update_start_
      -- 
    access_T_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(60) & access_T_CP_0_elements(285) & access_T_CP_0_elements(291) & access_T_CP_0_elements(299) & access_T_CP_0_elements(365);
      gj_access_T_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	32 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_sample_start__ps
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(32);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	33 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	34 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_update_start__ps
      -- 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(34);
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	35 
    -- CP-element group 60: 	283 
    -- CP-element group 60: 	289 
    -- CP-element group 60: 	297 
    -- CP-element group 60: 	364 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	56 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	28 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_loopback_trigger
      -- 
    access_T_CP_0_elements(61) <= access_T_CP_0_elements(28);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_loopback_sample_req_ps
      -- 
    phi_stmt_107_loopback_sample_req_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_107_loopback_sample_req_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => phi_stmt_107_req_1); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	29 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_entry_trigger
      -- 
    access_T_CP_0_elements(63) <= access_T_CP_0_elements(29);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_entry_sample_req_ps
      -- 
    phi_stmt_107_entry_sample_req_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_107_entry_sample_req_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(64), ack => phi_stmt_107_req_0); -- 
    -- Element group access_T_CP_0_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_phi_mux_ack_ps
      -- 
    phi_stmt_107_phi_mux_ack_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_107_ack_0, ack => access_T_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Sample/rr
      -- 
    rr_445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(68), ack => type_cast_110_inst_req_0); -- 
    access_T_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(66) & access_T_CP_0_elements(70);
      gj_access_T_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_update_start_
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Update/cr
      -- 
    cr_450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(69), ack => type_cast_110_inst_req_1); -- 
    access_T_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(67) & access_T_CP_0_elements(71);
      gj_access_T_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Sample/ra
      -- 
    ra_446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_110_inst_ack_0, ack => access_T_CP_0_elements(70)); -- 
    -- CP-element group 71:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_update_completed__ps
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Update/ca
      -- 
    ca_451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_110_inst_ack_1, ack => access_T_CP_0_elements(71)); -- 
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_sample_start__ps
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Sample/req
      -- 
    req_463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(72), ack => n_address2_308_111_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_update_start__ps
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_update_start_
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Update/req
      -- 
    req_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(73), ack => n_address2_308_111_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Sample/ack
      -- 
    ack_464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_308_111_buf_ack_0, ack => access_T_CP_0_elements(74)); -- 
    -- CP-element group 75:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Update/ack
      -- 
    ack_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_308_111_buf_ack_1, ack => access_T_CP_0_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	30 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	33 
    -- CP-element group 76: 	308 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	32 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_sample_start_
      -- 
    access_T_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(308);
      gj_access_T_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	30 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	81 
    -- CP-element group 77: 	313 
    -- CP-element group 77: 	319 
    -- CP-element group 77: 	327 
    -- CP-element group 77: 	368 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	34 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_update_start_
      -- 
    access_T_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(81) & access_T_CP_0_elements(313) & access_T_CP_0_elements(319) & access_T_CP_0_elements(327) & access_T_CP_0_elements(368);
      gj_access_T_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	32 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_sample_start__ps
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(32);
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	33 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	34 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_update_start__ps
      -- 
    access_T_CP_0_elements(80) <= access_T_CP_0_elements(34);
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	35 
    -- CP-element group 81: 	311 
    -- CP-element group 81: 	317 
    -- CP-element group 81: 	325 
    -- CP-element group 81: 	367 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	77 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	28 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_loopback_trigger
      -- 
    access_T_CP_0_elements(82) <= access_T_CP_0_elements(28);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_loopback_sample_req
      -- CP-element group 83: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_loopback_sample_req_ps
      -- 
    phi_stmt_112_loopback_sample_req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_112_loopback_sample_req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(83), ack => phi_stmt_112_req_1); -- 
    -- Element group access_T_CP_0_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	29 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_entry_trigger
      -- 
    access_T_CP_0_elements(84) <= access_T_CP_0_elements(29);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_entry_sample_req
      -- CP-element group 85: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_entry_sample_req_ps
      -- 
    phi_stmt_112_entry_sample_req_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_112_entry_sample_req_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(85), ack => phi_stmt_112_req_0); -- 
    -- Element group access_T_CP_0_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_phi_mux_ack
      -- CP-element group 86: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_phi_mux_ack_ps
      -- 
    phi_stmt_112_phi_mux_ack_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_112_ack_0, ack => access_T_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Sample/rr
      -- 
    rr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(89), ack => type_cast_115_inst_req_0); -- 
    access_T_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(87) & access_T_CP_0_elements(91);
      gj_access_T_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_update_start_
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Update/cr
      -- 
    cr_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(90), ack => type_cast_115_inst_req_1); -- 
    access_T_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(88) & access_T_CP_0_elements(92);
      gj_access_T_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_sample_completed__ps
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Sample/ra
      -- 
    ra_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_115_inst_ack_0, ack => access_T_CP_0_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_update_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Update/ca
      -- 
    ca_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_115_inst_ack_1, ack => access_T_CP_0_elements(92)); -- 
    -- CP-element group 93:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_sample_start__ps
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Sample/req
      -- 
    req_517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(93), ack => n_address3_380_116_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_update_start__ps
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_update_start_
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Update/req
      -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(94), ack => n_address3_380_116_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Sample/ack
      -- 
    ack_518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_380_116_buf_ack_0, ack => access_T_CP_0_elements(95)); -- 
    -- CP-element group 96:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Update/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_380_116_buf_ack_1, ack => access_T_CP_0_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	30 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	33 
    -- CP-element group 97: 	336 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	32 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_sample_start_
      -- 
    access_T_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(336);
      gj_access_T_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	30 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	102 
    -- CP-element group 98: 	341 
    -- CP-element group 98: 	347 
    -- CP-element group 98: 	355 
    -- CP-element group 98: 	371 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	34 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_update_start_
      -- 
    access_T_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(102) & access_T_CP_0_elements(341) & access_T_CP_0_elements(347) & access_T_CP_0_elements(355) & access_T_CP_0_elements(371);
      gj_access_T_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	32 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_sample_start__ps
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(32);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	33 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	34 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_update_start__ps
      -- 
    access_T_CP_0_elements(101) <= access_T_CP_0_elements(34);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	35 
    -- CP-element group 102: 	339 
    -- CP-element group 102: 	345 
    -- CP-element group 102: 	353 
    -- CP-element group 102: 	370 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	98 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	28 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_loopback_trigger
      -- 
    access_T_CP_0_elements(103) <= access_T_CP_0_elements(28);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_loopback_sample_req
      -- CP-element group 104: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_loopback_sample_req_ps
      -- 
    phi_stmt_117_loopback_sample_req_534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_117_loopback_sample_req_534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(104), ack => phi_stmt_117_req_1); -- 
    -- Element group access_T_CP_0_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	29 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_entry_trigger
      -- 
    access_T_CP_0_elements(105) <= access_T_CP_0_elements(29);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_entry_sample_req
      -- CP-element group 106: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_entry_sample_req_ps
      -- 
    phi_stmt_117_entry_sample_req_537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_117_entry_sample_req_537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(106), ack => phi_stmt_117_req_0); -- 
    -- Element group access_T_CP_0_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_phi_mux_ack
      -- CP-element group 107: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_phi_mux_ack_ps
      -- 
    phi_stmt_117_phi_mux_ack_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_117_ack_0, ack => access_T_CP_0_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Sample/rr
      -- 
    rr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(110), ack => type_cast_122_inst_req_0); -- 
    access_T_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(108) & access_T_CP_0_elements(112);
      gj_access_T_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_update_start_
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Update/cr
      -- 
    cr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(111), ack => type_cast_122_inst_req_1); -- 
    access_T_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(109) & access_T_CP_0_elements(113);
      gj_access_T_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_sample_completed__ps
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Sample/ra
      -- 
    ra_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_122_inst_ack_0, ack => access_T_CP_0_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_update_completed__ps
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Update/ca
      -- 
    ca_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_122_inst_ack_1, ack => access_T_CP_0_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Sample/req
      -- 
    req_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(114), ack => n_address4_452_123_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_update_start_
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Update/req
      -- 
    req_576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(115), ack => n_address4_452_123_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (4) 
      -- CP-element group 116: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_sample_completed__ps
      -- CP-element group 116: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Sample/ack
      -- 
    ack_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address4_452_123_buf_ack_0, ack => access_T_CP_0_elements(116)); -- 
    -- CP-element group 117:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_update_completed__ps
      -- CP-element group 117: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Update/ack
      -- 
    ack_577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address4_452_123_buf_ack_1, ack => access_T_CP_0_elements(117)); -- 
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	30 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	33 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	32 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_sample_start_
      -- 
    access_T_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33);
      gj_access_T_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	30 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	257 
    -- CP-element group 119: 	263 
    -- CP-element group 119: 	271 
    -- CP-element group 119: 	285 
    -- CP-element group 119: 	291 
    -- CP-element group 119: 	299 
    -- CP-element group 119: 	313 
    -- CP-element group 119: 	319 
    -- CP-element group 119: 	327 
    -- CP-element group 119: 	341 
    -- CP-element group 119: 	347 
    -- CP-element group 119: 	355 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	34 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_update_start_
      -- 
    access_T_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 1,6 => 0,7 => 0,8 => 1,9 => 0,10 => 0,11 => 1,12 => 0,13 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(123) & access_T_CP_0_elements(257) & access_T_CP_0_elements(263) & access_T_CP_0_elements(271) & access_T_CP_0_elements(285) & access_T_CP_0_elements(291) & access_T_CP_0_elements(299) & access_T_CP_0_elements(313) & access_T_CP_0_elements(319) & access_T_CP_0_elements(327) & access_T_CP_0_elements(341) & access_T_CP_0_elements(347) & access_T_CP_0_elements(355);
      gj_access_T_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	32 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_sample_start__ps
      -- 
    access_T_CP_0_elements(120) <= access_T_CP_0_elements(32);
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	33 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	34 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_update_start__ps
      -- 
    access_T_CP_0_elements(122) <= access_T_CP_0_elements(34);
    -- CP-element group 123:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	35 
    -- CP-element group 123: 	31 
    -- CP-element group 123: 	255 
    -- CP-element group 123: 	261 
    -- CP-element group 123: 	269 
    -- CP-element group 123: 	283 
    -- CP-element group 123: 	289 
    -- CP-element group 123: 	297 
    -- CP-element group 123: 	311 
    -- CP-element group 123: 	317 
    -- CP-element group 123: 	325 
    -- CP-element group 123: 	339 
    -- CP-element group 123: 	345 
    -- CP-element group 123: 	353 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	119 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	28 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_loopback_trigger
      -- 
    access_T_CP_0_elements(124) <= access_T_CP_0_elements(28);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_loopback_sample_req
      -- CP-element group 125: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_loopback_sample_req_ps
      -- 
    phi_stmt_124_loopback_sample_req_588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_124_loopback_sample_req_588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(125), ack => phi_stmt_124_req_1); -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	29 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_entry_trigger
      -- 
    access_T_CP_0_elements(126) <= access_T_CP_0_elements(29);
    -- CP-element group 127:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_entry_sample_req
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_entry_sample_req_ps
      -- 
    phi_stmt_124_entry_sample_req_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_124_entry_sample_req_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(127), ack => phi_stmt_124_req_0); -- 
    -- Element group access_T_CP_0_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_phi_mux_ack
      -- CP-element group 128: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_phi_mux_ack_ps
      -- 
    phi_stmt_124_phi_mux_ack_594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_124_ack_0, ack => access_T_CP_0_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (4) 
      -- CP-element group 129: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_sample_start__ps
      -- CP-element group 129: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_sample_completed__ps
      -- CP-element group 129: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_update_start__ps
      -- CP-element group 130: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_update_start_
      -- 
    -- Element group access_T_CP_0_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_update_completed__ps
      -- 
    access_T_CP_0_elements(131) <= access_T_CP_0_elements(132);
    -- CP-element group 132:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	131 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(132) is a control-delay.
    cp_element_132_delay: control_delay_element  generic map(name => " 132_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(130), ack => access_T_CP_0_elements(132), clk => clk, reset =>reset);
    -- CP-element group 133:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Sample/req
      -- 
    req_615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(133), ack => n_mycounter_168_128_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_update_start__ps
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_update_start_
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Update/req
      -- 
    req_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(134), ack => n_mycounter_168_128_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (4) 
      -- CP-element group 135: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_sample_completed__ps
      -- CP-element group 135: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Sample/ack
      -- 
    ack_616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter_168_128_buf_ack_0, ack => access_T_CP_0_elements(135)); -- 
    -- CP-element group 136:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (4) 
      -- CP-element group 136: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_update_completed__ps
      -- CP-element group 136: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Update/ack
      -- 
    ack_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter_168_128_buf_ack_1, ack => access_T_CP_0_elements(136)); -- 
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	30 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	33 
    -- CP-element group 137: 	268 
    -- CP-element group 137: 	272 
    -- CP-element group 137: 	276 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	32 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_sample_start_
      -- 
    access_T_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(268) & access_T_CP_0_elements(272) & access_T_CP_0_elements(276);
      gj_access_T_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	30 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: 	275 
    -- CP-element group 138: 	362 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	34 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_update_start_
      -- 
    access_T_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(140) & access_T_CP_0_elements(275) & access_T_CP_0_elements(362);
      gj_access_T_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	33 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(139) is bound as output of CP function.
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	35 
    -- CP-element group 140: 	273 
    -- CP-element group 140: 	361 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	138 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	28 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_loopback_trigger
      -- 
    access_T_CP_0_elements(141) <= access_T_CP_0_elements(28);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_loopback_sample_req_ps
      -- 
    phi_stmt_129_loopback_sample_req_632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_129_loopback_sample_req_632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(142), ack => phi_stmt_129_req_1); -- 
    -- Element group access_T_CP_0_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	29 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_entry_trigger
      -- 
    access_T_CP_0_elements(143) <= access_T_CP_0_elements(29);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_entry_sample_req_ps
      -- 
    phi_stmt_129_entry_sample_req_635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_129_entry_sample_req_635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(144), ack => phi_stmt_129_req_0); -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_phi_mux_ack_ps
      -- 
    phi_stmt_129_phi_mux_ack_638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_129_ack_0, ack => access_T_CP_0_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Sample/req
      -- 
    req_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(146), ack => my_fetch1_53_131_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (4) 
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_update_start_
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Update/req
      -- 
    req_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(147), ack => my_fetch1_53_131_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (4) 
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_sample_completed__ps
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Sample/ack
      -- 
    ack_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch1_53_131_buf_ack_0, ack => access_T_CP_0_elements(148)); -- 
    -- CP-element group 149:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (4) 
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_update_completed__ps
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Update/ack
      -- 
    ack_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch1_53_131_buf_ack_1, ack => access_T_CP_0_elements(149)); -- 
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_sample_start_
      -- 
    req_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => n_fetch_val1_276_132_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Update/req
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_update_start_
      -- 
    req_674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(151), ack => n_fetch_val1_276_132_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Sample/ack
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_sample_completed_
      -- 
    ack_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val1_276_132_buf_ack_0, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Update/ack
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_update_completed__ps
      -- 
    ack_675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val1_276_132_buf_ack_1, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  join  transition  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	30 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	33 
    -- CP-element group 154: 	296 
    -- CP-element group 154: 	300 
    -- CP-element group 154: 	304 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	32 
    -- CP-element group 154:  members (1) 
      -- CP-element group 154: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_sample_start_
      -- 
    access_T_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(296) & access_T_CP_0_elements(300) & access_T_CP_0_elements(304);
      gj_access_T_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	30 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	159 
    -- CP-element group 155: 	303 
    -- CP-element group 155: 	365 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	34 
    -- CP-element group 155:  members (1) 
      -- CP-element group 155: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_update_start_
      -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(159) & access_T_CP_0_elements(303) & access_T_CP_0_elements(365);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	32 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (1) 
      -- CP-element group 156: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_sample_start__ps
      -- 
    access_T_CP_0_elements(156) <= access_T_CP_0_elements(32);
    -- CP-element group 157:  join  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	33 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(157) is bound as output of CP function.
    -- CP-element group 158:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	34 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_update_start__ps
      -- 
    access_T_CP_0_elements(158) <= access_T_CP_0_elements(34);
    -- CP-element group 159:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	35 
    -- CP-element group 159: 	301 
    -- CP-element group 159: 	364 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	155 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(159) is bound as output of CP function.
    -- CP-element group 160:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	28 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_loopback_trigger
      -- 
    access_T_CP_0_elements(160) <= access_T_CP_0_elements(28);
    -- CP-element group 161:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (2) 
      -- CP-element group 161: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_loopback_sample_req
      -- CP-element group 161: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_loopback_sample_req_ps
      -- 
    phi_stmt_133_loopback_sample_req_686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_133_loopback_sample_req_686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(161), ack => phi_stmt_133_req_1); -- 
    -- Element group access_T_CP_0_elements(161) is bound as output of CP function.
    -- CP-element group 162:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	29 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_entry_trigger
      -- 
    access_T_CP_0_elements(162) <= access_T_CP_0_elements(29);
    -- CP-element group 163:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_entry_sample_req
      -- CP-element group 163: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_entry_sample_req_ps
      -- 
    phi_stmt_133_entry_sample_req_689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_133_entry_sample_req_689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => phi_stmt_133_req_0); -- 
    -- Element group access_T_CP_0_elements(163) is bound as output of CP function.
    -- CP-element group 164:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_phi_mux_ack
      -- CP-element group 164: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_phi_mux_ack_ps
      -- 
    phi_stmt_133_phi_mux_ack_692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_133_ack_0, ack => access_T_CP_0_elements(164)); -- 
    -- CP-element group 165:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (4) 
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_sample_start__ps
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Sample/req
      -- 
    req_705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(165), ack => my_fetch2_67_135_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(165) is bound as output of CP function.
    -- CP-element group 166:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (4) 
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_update_start__ps
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_update_start_
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Update/req
      -- 
    req_710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(166), ack => my_fetch2_67_135_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(166) is bound as output of CP function.
    -- CP-element group 167:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (4) 
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_sample_completed__ps
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Sample/ack
      -- 
    ack_706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch2_67_135_buf_ack_0, ack => access_T_CP_0_elements(167)); -- 
    -- CP-element group 168:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (4) 
      -- CP-element group 168: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_update_completed__ps
      -- CP-element group 168: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Update/ack
      -- 
    ack_711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch2_67_135_buf_ack_1, ack => access_T_CP_0_elements(168)); -- 
    -- CP-element group 169:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (4) 
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_sample_start__ps
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Sample/req
      -- 
    req_723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(169), ack => n_fetch_val2_348_136_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(169) is bound as output of CP function.
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_update_start__ps
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_update_start_
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Update/req
      -- 
    req_728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(170), ack => n_fetch_val2_348_136_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(170) is bound as output of CP function.
    -- CP-element group 171:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (4) 
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_sample_completed__ps
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Sample/ack
      -- 
    ack_724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val2_348_136_buf_ack_0, ack => access_T_CP_0_elements(171)); -- 
    -- CP-element group 172:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (4) 
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_update_completed__ps
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Update/ack
      -- 
    ack_729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val2_348_136_buf_ack_1, ack => access_T_CP_0_elements(172)); -- 
    -- CP-element group 173:  join  transition  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	30 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	33 
    -- CP-element group 173: 	324 
    -- CP-element group 173: 	328 
    -- CP-element group 173: 	332 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	32 
    -- CP-element group 173:  members (1) 
      -- CP-element group 173: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_sample_start_
      -- 
    access_T_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(324) & access_T_CP_0_elements(328) & access_T_CP_0_elements(332);
      gj_access_T_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	30 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	178 
    -- CP-element group 174: 	331 
    -- CP-element group 174: 	368 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	34 
    -- CP-element group 174:  members (1) 
      -- CP-element group 174: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_update_start_
      -- 
    access_T_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(178) & access_T_CP_0_elements(331) & access_T_CP_0_elements(368);
      gj_access_T_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	32 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_sample_start__ps
      -- 
    access_T_CP_0_elements(175) <= access_T_CP_0_elements(32);
    -- CP-element group 176:  join  transition  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	33 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(176) is bound as output of CP function.
    -- CP-element group 177:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	34 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_update_start__ps
      -- 
    access_T_CP_0_elements(177) <= access_T_CP_0_elements(34);
    -- CP-element group 178:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	35 
    -- CP-element group 178: 	329 
    -- CP-element group 178: 	367 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	174 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(178) is bound as output of CP function.
    -- CP-element group 179:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	28 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_loopback_trigger
      -- 
    access_T_CP_0_elements(179) <= access_T_CP_0_elements(28);
    -- CP-element group 180:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_loopback_sample_req
      -- CP-element group 180: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_loopback_sample_req_ps
      -- 
    phi_stmt_137_loopback_sample_req_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_137_loopback_sample_req_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => phi_stmt_137_req_1); -- 
    -- Element group access_T_CP_0_elements(180) is bound as output of CP function.
    -- CP-element group 181:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	29 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_entry_trigger
      -- 
    access_T_CP_0_elements(181) <= access_T_CP_0_elements(29);
    -- CP-element group 182:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (2) 
      -- CP-element group 182: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_entry_sample_req
      -- CP-element group 182: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_entry_sample_req_ps
      -- 
    phi_stmt_137_entry_sample_req_743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_137_entry_sample_req_743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => phi_stmt_137_req_0); -- 
    -- Element group access_T_CP_0_elements(182) is bound as output of CP function.
    -- CP-element group 183:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_phi_mux_ack
      -- CP-element group 183: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_phi_mux_ack_ps
      -- 
    phi_stmt_137_phi_mux_ack_746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_137_ack_0, ack => access_T_CP_0_elements(183)); -- 
    -- CP-element group 184:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (4) 
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_sample_start__ps
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Sample/req
      -- 
    req_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(184), ack => my_fetch3_81_139_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(184) is bound as output of CP function.
    -- CP-element group 185:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (4) 
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_update_start__ps
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_update_start_
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Update/req
      -- 
    req_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(185), ack => my_fetch3_81_139_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(185) is bound as output of CP function.
    -- CP-element group 186:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (4) 
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_sample_completed__ps
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Sample/ack
      -- 
    ack_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch3_81_139_buf_ack_0, ack => access_T_CP_0_elements(186)); -- 
    -- CP-element group 187:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (4) 
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_update_completed__ps
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Update/ack
      -- 
    ack_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch3_81_139_buf_ack_1, ack => access_T_CP_0_elements(187)); -- 
    -- CP-element group 188:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (4) 
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_sample_start__ps
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Sample/req
      -- 
    req_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(188), ack => n_fetch_val3_420_140_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(188) is bound as output of CP function.
    -- CP-element group 189:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (4) 
      -- CP-element group 189: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_update_start__ps
      -- CP-element group 189: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_update_start_
      -- CP-element group 189: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Update/req
      -- 
    req_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(189), ack => n_fetch_val3_420_140_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(189) is bound as output of CP function.
    -- CP-element group 190:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (4) 
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_sample_completed__ps
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Sample/ack
      -- 
    ack_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val3_420_140_buf_ack_0, ack => access_T_CP_0_elements(190)); -- 
    -- CP-element group 191:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (4) 
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_update_completed__ps
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Update/ack
      -- 
    ack_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val3_420_140_buf_ack_1, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  join  transition  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	30 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	33 
    -- CP-element group 192: 	352 
    -- CP-element group 192: 	356 
    -- CP-element group 192: 	360 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	32 
    -- CP-element group 192:  members (1) 
      -- CP-element group 192: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_sample_start_
      -- 
    access_T_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(352) & access_T_CP_0_elements(356) & access_T_CP_0_elements(360);
      gj_access_T_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	30 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	197 
    -- CP-element group 193: 	359 
    -- CP-element group 193: 	371 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	34 
    -- CP-element group 193:  members (1) 
      -- CP-element group 193: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_update_start_
      -- 
    access_T_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(197) & access_T_CP_0_elements(359) & access_T_CP_0_elements(371);
      gj_access_T_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	32 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (1) 
      -- CP-element group 194: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_sample_start__ps
      -- 
    access_T_CP_0_elements(194) <= access_T_CP_0_elements(32);
    -- CP-element group 195:  join  transition  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	33 
    -- CP-element group 195:  members (1) 
      -- CP-element group 195: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(195) is bound as output of CP function.
    -- CP-element group 196:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	34 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (1) 
      -- CP-element group 196: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_update_start__ps
      -- 
    access_T_CP_0_elements(196) <= access_T_CP_0_elements(34);
    -- CP-element group 197:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	35 
    -- CP-element group 197: 	357 
    -- CP-element group 197: 	370 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	193 
    -- CP-element group 197:  members (2) 
      -- CP-element group 197: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(197) is bound as output of CP function.
    -- CP-element group 198:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	28 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_loopback_trigger
      -- 
    access_T_CP_0_elements(198) <= access_T_CP_0_elements(28);
    -- CP-element group 199:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_loopback_sample_req
      -- CP-element group 199: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_loopback_sample_req_ps
      -- 
    phi_stmt_141_loopback_sample_req_794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_141_loopback_sample_req_794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(199), ack => phi_stmt_141_req_1); -- 
    -- Element group access_T_CP_0_elements(199) is bound as output of CP function.
    -- CP-element group 200:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	29 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_entry_trigger
      -- 
    access_T_CP_0_elements(200) <= access_T_CP_0_elements(29);
    -- CP-element group 201:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (2) 
      -- CP-element group 201: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_entry_sample_req
      -- CP-element group 201: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_entry_sample_req_ps
      -- 
    phi_stmt_141_entry_sample_req_797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_141_entry_sample_req_797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => phi_stmt_141_req_0); -- 
    -- Element group access_T_CP_0_elements(201) is bound as output of CP function.
    -- CP-element group 202:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (2) 
      -- CP-element group 202: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_phi_mux_ack
      -- CP-element group 202: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_phi_mux_ack_ps
      -- 
    phi_stmt_141_phi_mux_ack_800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_141_ack_0, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (4) 
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_sample_start__ps
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Sample/req
      -- 
    req_813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(203), ack => my_fetch4_99_143_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(203) is bound as output of CP function.
    -- CP-element group 204:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (4) 
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_update_start__ps
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_update_start_
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Update/req
      -- 
    req_818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(204), ack => my_fetch4_99_143_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(204) is bound as output of CP function.
    -- CP-element group 205:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (4) 
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_sample_completed__ps
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Sample/ack
      -- 
    ack_814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch4_99_143_buf_ack_0, ack => access_T_CP_0_elements(205)); -- 
    -- CP-element group 206:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (4) 
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_update_completed__ps
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Update/ack
      -- 
    ack_819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch4_99_143_buf_ack_1, ack => access_T_CP_0_elements(206)); -- 
    -- CP-element group 207:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (4) 
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_sample_start__ps
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Sample/req
      -- 
    req_831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(207), ack => n_fetch_val4_492_144_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(207) is bound as output of CP function.
    -- CP-element group 208:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (4) 
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_update_start__ps
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_update_start_
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Update/req
      -- 
    req_836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(208), ack => n_fetch_val4_492_144_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(208) is bound as output of CP function.
    -- CP-element group 209:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (4) 
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_sample_completed__ps
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Sample/ack
      -- 
    ack_832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val4_492_144_buf_ack_0, ack => access_T_CP_0_elements(209)); -- 
    -- CP-element group 210:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (4) 
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_update_completed__ps
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Update/ack
      -- 
    ack_837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val4_492_144_buf_ack_1, ack => access_T_CP_0_elements(210)); -- 
    -- CP-element group 211:  join  transition  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	30 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	33 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	32 
    -- CP-element group 211:  members (1) 
      -- CP-element group 211: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_sample_start_
      -- 
    access_T_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33);
      gj_access_T_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  join  transition  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	30 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	216 
    -- CP-element group 212: 	263 
    -- CP-element group 212: 	271 
    -- CP-element group 212: 	291 
    -- CP-element group 212: 	299 
    -- CP-element group 212: 	319 
    -- CP-element group 212: 	327 
    -- CP-element group 212: 	362 
    -- CP-element group 212: 	365 
    -- CP-element group 212: 	368 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	34 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_update_start_
      -- 
    access_T_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(216) & access_T_CP_0_elements(263) & access_T_CP_0_elements(271) & access_T_CP_0_elements(291) & access_T_CP_0_elements(299) & access_T_CP_0_elements(319) & access_T_CP_0_elements(327) & access_T_CP_0_elements(362) & access_T_CP_0_elements(365) & access_T_CP_0_elements(368);
      gj_access_T_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	32 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_sample_start__ps
      -- 
    access_T_CP_0_elements(213) <= access_T_CP_0_elements(32);
    -- CP-element group 214:  join  transition  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	33 
    -- CP-element group 214:  members (1) 
      -- CP-element group 214: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(214) is bound as output of CP function.
    -- CP-element group 215:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	34 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_update_start__ps
      -- 
    access_T_CP_0_elements(215) <= access_T_CP_0_elements(34);
    -- CP-element group 216:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	35 
    -- CP-element group 216: 	31 
    -- CP-element group 216: 	261 
    -- CP-element group 216: 	269 
    -- CP-element group 216: 	289 
    -- CP-element group 216: 	297 
    -- CP-element group 216: 	317 
    -- CP-element group 216: 	325 
    -- CP-element group 216: 	361 
    -- CP-element group 216: 	364 
    -- CP-element group 216: 	367 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	212 
    -- CP-element group 216:  members (2) 
      -- CP-element group 216: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(216) is bound as output of CP function.
    -- CP-element group 217:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	28 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (1) 
      -- CP-element group 217: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_loopback_trigger
      -- 
    access_T_CP_0_elements(217) <= access_T_CP_0_elements(28);
    -- CP-element group 218:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_loopback_sample_req
      -- CP-element group 218: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_loopback_sample_req_ps
      -- 
    phi_stmt_145_loopback_sample_req_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_145_loopback_sample_req_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(218), ack => phi_stmt_145_req_1); -- 
    -- Element group access_T_CP_0_elements(218) is bound as output of CP function.
    -- CP-element group 219:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	29 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (1) 
      -- CP-element group 219: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_entry_trigger
      -- 
    access_T_CP_0_elements(219) <= access_T_CP_0_elements(29);
    -- CP-element group 220:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (2) 
      -- CP-element group 220: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_entry_sample_req
      -- CP-element group 220: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_entry_sample_req_ps
      -- 
    phi_stmt_145_entry_sample_req_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_145_entry_sample_req_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(220), ack => phi_stmt_145_req_0); -- 
    -- Element group access_T_CP_0_elements(220) is bound as output of CP function.
    -- CP-element group 221:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (2) 
      -- CP-element group 221: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_phi_mux_ack
      -- CP-element group 221: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_phi_mux_ack_ps
      -- 
    phi_stmt_145_phi_mux_ack_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_145_ack_0, ack => access_T_CP_0_elements(221)); -- 
    -- CP-element group 222:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (4) 
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_sample_start__ps
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_sample_completed__ps
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(222) is bound as output of CP function.
    -- CP-element group 223:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (2) 
      -- CP-element group 223: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_update_start__ps
      -- CP-element group 223: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_update_start_
      -- 
    -- Element group access_T_CP_0_elements(223) is bound as output of CP function.
    -- CP-element group 224:  join  transition  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	225 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (1) 
      -- CP-element group 224: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_update_completed__ps
      -- 
    access_T_CP_0_elements(224) <= access_T_CP_0_elements(225);
    -- CP-element group 225:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	224 
    -- CP-element group 225:  members (1) 
      -- CP-element group 225: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(225) is a control-delay.
    cp_element_225_delay: control_delay_element  generic map(name => " 225_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(223), ack => access_T_CP_0_elements(225), clk => clk, reset =>reset);
    -- CP-element group 226:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (4) 
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_sample_start__ps
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Sample/req
      -- 
    req_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(226), ack => n_row1_186_149_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(226) is bound as output of CP function.
    -- CP-element group 227:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (4) 
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_update_start__ps
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_update_start_
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Update/req
      -- 
    req_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(227), ack => n_row1_186_149_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(227) is bound as output of CP function.
    -- CP-element group 228:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (4) 
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_sample_completed__ps
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Sample/ack
      -- 
    ack_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_186_149_buf_ack_0, ack => access_T_CP_0_elements(228)); -- 
    -- CP-element group 229:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (4) 
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_update_completed__ps
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Update/ack
      -- 
    ack_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_186_149_buf_ack_1, ack => access_T_CP_0_elements(229)); -- 
    -- CP-element group 230:  join  transition  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	30 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	33 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	32 
    -- CP-element group 230:  members (1) 
      -- CP-element group 230: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_sample_start_
      -- 
    access_T_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33);
      gj_access_T_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	30 
    -- CP-element group 231: marked-predecessors 
    -- CP-element group 231: 	235 
    -- CP-element group 231: 	347 
    -- CP-element group 231: 	355 
    -- CP-element group 231: 	371 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	34 
    -- CP-element group 231:  members (1) 
      -- CP-element group 231: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_update_start_
      -- 
    access_T_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(235) & access_T_CP_0_elements(347) & access_T_CP_0_elements(355) & access_T_CP_0_elements(371);
      gj_access_T_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	32 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_sample_start__ps
      -- 
    access_T_CP_0_elements(232) <= access_T_CP_0_elements(32);
    -- CP-element group 233:  join  transition  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	33 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(233) is bound as output of CP function.
    -- CP-element group 234:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	34 
    -- CP-element group 234: successors 
    -- CP-element group 234:  members (1) 
      -- CP-element group 234: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_update_start__ps
      -- 
    access_T_CP_0_elements(234) <= access_T_CP_0_elements(34);
    -- CP-element group 235:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	35 
    -- CP-element group 235: 	345 
    -- CP-element group 235: 	353 
    -- CP-element group 235: 	370 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	231 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(235) is bound as output of CP function.
    -- CP-element group 236:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	28 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_loopback_trigger
      -- 
    access_T_CP_0_elements(236) <= access_T_CP_0_elements(28);
    -- CP-element group 237:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (2) 
      -- CP-element group 237: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_loopback_sample_req
      -- CP-element group 237: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_loopback_sample_req_ps
      -- 
    phi_stmt_150_loopback_sample_req_892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_150_loopback_sample_req_892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(237), ack => phi_stmt_150_req_1); -- 
    -- Element group access_T_CP_0_elements(237) is bound as output of CP function.
    -- CP-element group 238:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	29 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (1) 
      -- CP-element group 238: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_entry_trigger
      -- 
    access_T_CP_0_elements(238) <= access_T_CP_0_elements(29);
    -- CP-element group 239:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_entry_sample_req
      -- CP-element group 239: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_entry_sample_req_ps
      -- 
    phi_stmt_150_entry_sample_req_895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_150_entry_sample_req_895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(239), ack => phi_stmt_150_req_0); -- 
    -- Element group access_T_CP_0_elements(239) is bound as output of CP function.
    -- CP-element group 240:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_phi_mux_ack
      -- CP-element group 240: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_phi_mux_ack_ps
      -- 
    phi_stmt_150_phi_mux_ack_898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_150_ack_0, ack => access_T_CP_0_elements(240)); -- 
    -- CP-element group 241:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (4) 
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_sample_start__ps
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_sample_completed__ps
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(241) is bound as output of CP function.
    -- CP-element group 242:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_update_start__ps
      -- CP-element group 242: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_update_start_
      -- 
    -- Element group access_T_CP_0_elements(242) is bound as output of CP function.
    -- CP-element group 243:  join  transition  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	244 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (1) 
      -- CP-element group 243: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_update_completed__ps
      -- 
    access_T_CP_0_elements(243) <= access_T_CP_0_elements(244);
    -- CP-element group 244:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	243 
    -- CP-element group 244:  members (1) 
      -- CP-element group 244: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(244) is a control-delay.
    cp_element_244_delay: control_delay_element  generic map(name => " 244_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(242), ack => access_T_CP_0_elements(244), clk => clk, reset =>reset);
    -- CP-element group 245:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (4) 
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_sample_start__ps
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Sample/req
      -- 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(245), ack => n_row2_194_154_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(245) is bound as output of CP function.
    -- CP-element group 246:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (4) 
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_update_start__ps
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_update_start_
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Update/req
      -- 
    req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(246), ack => n_row2_194_154_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(246) is bound as output of CP function.
    -- CP-element group 247:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (4) 
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_sample_completed__ps
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Sample/ack
      -- 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_194_154_buf_ack_0, ack => access_T_CP_0_elements(247)); -- 
    -- CP-element group 248:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (4) 
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_update_completed__ps
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Update/ack
      -- 
    ack_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_194_154_buf_ack_1, ack => access_T_CP_0_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	30 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Sample/rr
      -- 
    rr_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(249), ack => type_cast_227_inst_req_0); -- 
    access_T_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(251);
      gj_access_T_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	33 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	252 
    -- CP-element group 250: 	257 
    -- CP-element group 250: 	263 
    -- CP-element group 250: 	271 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_update_start_
      -- CP-element group 250: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Update/cr
      -- 
    cr_939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(250), ack => type_cast_227_inst_req_1); -- 
    access_T_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(252) & access_T_CP_0_elements(257) & access_T_CP_0_elements(263) & access_T_CP_0_elements(271);
      gj_access_T_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Sample/ra
      -- 
    ra_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_227_inst_ack_0, ack => access_T_CP_0_elements(251)); -- 
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	255 
    -- CP-element group 252: 	261 
    -- CP-element group 252: 	269 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	36 
    -- CP-element group 252: 	250 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Update/ca
      -- 
    ca_940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_227_inst_ack_1, ack => access_T_CP_0_elements(252)); -- 
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	258 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	259 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	259 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_request/req
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_request/$entry
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_sample_start_
      -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(253), ack => addr_of_255_final_reg_req_0); -- 
    access_T_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(258) & access_T_CP_0_elements(259);
      gj_access_T_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	30 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	260 
    -- CP-element group 254: 	267 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	260 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_complete/$entry
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_complete/req
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_update_start_
      -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(254), ack => addr_of_255_final_reg_req_1); -- 
    access_T_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(260) & access_T_CP_0_elements(267);
      gj_access_T_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	41 
    -- CP-element group 255: 	123 
    -- CP-element group 255: 	252 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (13) 
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_resized_1
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_scaled_1
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_computed_1
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_resize_1/$entry
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_resize_1/$exit
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_resize_1/index_resize_req
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_resize_1/index_resize_ack
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_scale_1/$entry
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_scale_1/$exit
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_scale_1/scale_rename_req
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_scale_1/scale_rename_ack
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Sample/req
      -- 
    req_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(255), ack => array_obj_ref_254_index_offset_req_0); -- 
    access_T_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(41) & access_T_CP_0_elements(123) & access_T_CP_0_elements(252);
      gj_access_T_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	30 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: 	259 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_update_start
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Update/req
      -- 
    req_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(256), ack => array_obj_ref_254_index_offset_req_1); -- 
    access_T_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(258) & access_T_CP_0_elements(259);
      gj_access_T_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	374 
    -- CP-element group 257: marked-successors 
    -- CP-element group 257: 	37 
    -- CP-element group 257: 	119 
    -- CP-element group 257: 	250 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_sample_complete
      -- CP-element group 257: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Sample/ack
      -- 
    ack_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_254_index_offset_ack_0, ack => access_T_CP_0_elements(257)); -- 
    -- CP-element group 258:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	253 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (8) 
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_base_plus_offset/sum_rename_ack
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_base_plus_offset/sum_rename_req
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_base_plus_offset/$exit
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_base_plus_offset/$entry
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_root_address_calculated
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_offset_calculated
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Update/ack
      -- 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_254_index_offset_ack_1, ack => access_T_CP_0_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	253 
    -- CP-element group 259: successors 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	253 
    -- CP-element group 259: 	256 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_request/ack
      -- CP-element group 259: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_request/$exit
      -- CP-element group 259: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_sample_completed_
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_255_final_reg_ack_0, ack => access_T_CP_0_elements(259)); -- 
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	254 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	265 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	254 
    -- CP-element group 260:  members (19) 
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_complete/$exit
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_word_addrgen/root_register_ack
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_word_addrgen/root_register_req
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_word_addrgen/$exit
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_word_addrgen/$entry
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_plus_offset/sum_rename_ack
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_complete/ack
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_plus_offset/sum_rename_req
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_plus_offset/$exit
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_plus_offset/$entry
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_addr_resize/base_resize_ack
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_addr_resize/base_resize_req
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_addr_resize/$exit
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_addr_resize/$entry
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_address_resized
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_root_address_calculated
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_word_address_calculated
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_address_calculated
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_update_completed_
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_255_final_reg_ack_1, ack => access_T_CP_0_elements(260)); -- 
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	41 
    -- CP-element group 261: 	123 
    -- CP-element group 261: 	216 
    -- CP-element group 261: 	252 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Sample/req
      -- CP-element group 261: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Sample/$entry
      -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(261), ack => W_fn1_254_delayed_7_0_257_inst_req_0); -- 
    access_T_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(41) & access_T_CP_0_elements(123) & access_T_CP_0_elements(216) & access_T_CP_0_elements(252) & access_T_CP_0_elements(263);
      gj_access_T_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	264 
    -- CP-element group 262: 	267 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_update_start_
      -- CP-element group 262: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Update/req
      -- CP-element group 262: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Update/$entry
      -- 
    req_999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(262), ack => W_fn1_254_delayed_7_0_257_inst_req_1); -- 
    access_T_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(264) & access_T_CP_0_elements(267);
      gj_access_T_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	37 
    -- CP-element group 263: 	119 
    -- CP-element group 263: 	212 
    -- CP-element group 263: 	250 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Sample/$exit
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_254_delayed_7_0_257_inst_ack_0, ack => access_T_CP_0_elements(263)); -- 
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_update_completed_
      -- 
    ack_1000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_254_delayed_7_0_257_inst_ack_1, ack => access_T_CP_0_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	260 
    -- CP-element group 265: 	264 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (5) 
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/word_0/rr
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/word_0/$entry
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/$entry
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_sample_start_
      -- 
    rr_1033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(265), ack => ptr_deref_263_load_0_req_0); -- 
    access_T_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(260) & access_T_CP_0_elements(264) & access_T_CP_0_elements(267);
      gj_access_T_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	33 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (5) 
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/word_0/cr
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/word_0/$entry
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/$entry
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_update_start_
      -- 
    cr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(266), ack => ptr_deref_263_load_0_req_1); -- 
    access_T_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(268);
      gj_access_T_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	254 
    -- CP-element group 267: 	262 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (5) 
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/word_0/ra
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/word_0/$exit
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/$exit
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_sample_completed_
      -- 
    ra_1034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_load_0_ack_0, ack => access_T_CP_0_elements(267)); -- 
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	374 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	137 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (9) 
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/ptr_deref_263_Merge/merge_req
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/ptr_deref_263_Merge/$exit
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/ptr_deref_263_Merge/$entry
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/word_0/ca
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/word_0/$exit
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/$exit
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/ptr_deref_263_Merge/merge_ack
      -- 
    ca_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_load_0_ack_1, ack => access_T_CP_0_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	41 
    -- CP-element group 269: 	123 
    -- CP-element group 269: 	216 
    -- CP-element group 269: 	252 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Sample/req
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_sample_start_
      -- 
    req_1058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(269), ack => W_fn1_260_delayed_13_0_265_inst_req_0); -- 
    access_T_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(41) & access_T_CP_0_elements(123) & access_T_CP_0_elements(216) & access_T_CP_0_elements(252) & access_T_CP_0_elements(271);
      gj_access_T_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	33 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	272 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Update/req
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_update_start_
      -- 
    req_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(270), ack => W_fn1_260_delayed_13_0_265_inst_req_1); -- 
    access_T_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(272);
      gj_access_T_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	37 
    -- CP-element group 271: 	119 
    -- CP-element group 271: 	212 
    -- CP-element group 271: 	250 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_sample_completed_
      -- 
    ack_1059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_260_delayed_13_0_265_inst_ack_0, ack => access_T_CP_0_elements(271)); -- 
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	374 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	137 
    -- CP-element group 272: 	270 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_update_completed_
      -- 
    ack_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_260_delayed_13_0_265_inst_ack_1, ack => access_T_CP_0_elements(272)); -- 
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	140 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Sample/req
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_sample_start_
      -- 
    req_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(273), ack => W_fetch_val1_262_delayed_13_0_268_inst_req_0); -- 
    access_T_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(140) & access_T_CP_0_elements(275);
      gj_access_T_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	33 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	276 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Update/req
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_update_start_
      -- 
    req_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(274), ack => W_fetch_val1_262_delayed_13_0_268_inst_req_1); -- 
    access_T_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(276);
      gj_access_T_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	138 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_sample_completed_
      -- 
    ack_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val1_262_delayed_13_0_268_inst_ack_0, ack => access_T_CP_0_elements(275)); -- 
    -- CP-element group 276:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	374 
    -- CP-element group 276: marked-successors 
    -- CP-element group 276: 	137 
    -- CP-element group 276: 	274 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_update_completed_
      -- 
    ack_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val1_262_delayed_13_0_268_inst_ack_1, ack => access_T_CP_0_elements(276)); -- 
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	30 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Sample/rr
      -- CP-element group 277: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_sample_start_
      -- 
    rr_1086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(277), ack => type_cast_299_inst_req_0); -- 
    access_T_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(279);
      gj_access_T_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	33 
    -- CP-element group 278: marked-predecessors 
    -- CP-element group 278: 	280 
    -- CP-element group 278: 	285 
    -- CP-element group 278: 	291 
    -- CP-element group 278: 	299 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Update/cr
      -- CP-element group 278: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Update/$entry
      -- CP-element group 278: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_update_start_
      -- 
    cr_1091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(278), ack => type_cast_299_inst_req_1); -- 
    access_T_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(280) & access_T_CP_0_elements(285) & access_T_CP_0_elements(291) & access_T_CP_0_elements(299);
      gj_access_T_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Sample/ra
      -- CP-element group 279: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_sample_completed_
      -- 
    ra_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_299_inst_ack_0, ack => access_T_CP_0_elements(279)); -- 
    -- CP-element group 280:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280: 	289 
    -- CP-element group 280: 	297 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	55 
    -- CP-element group 280: 	278 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Update/ca
      -- CP-element group 280: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_update_completed_
      -- 
    ca_1092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_299_inst_ack_1, ack => access_T_CP_0_elements(280)); -- 
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	286 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	287 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	287 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_request/req
      -- CP-element group 281: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_request/$entry
      -- CP-element group 281: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_sample_start_
      -- 
    req_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(281), ack => addr_of_327_final_reg_req_0); -- 
    access_T_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(286) & access_T_CP_0_elements(287);
      gj_access_T_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	30 
    -- CP-element group 282: marked-predecessors 
    -- CP-element group 282: 	288 
    -- CP-element group 282: 	295 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	288 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_complete/req
      -- CP-element group 282: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_complete/$entry
      -- CP-element group 282: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_update_start_
      -- 
    req_1137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(282), ack => addr_of_327_final_reg_req_1); -- 
    access_T_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(288) & access_T_CP_0_elements(295);
      gj_access_T_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	60 
    -- CP-element group 283: 	123 
    -- CP-element group 283: 	280 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	285 
    -- CP-element group 283:  members (13) 
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_scale_1/scale_rename_ack
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_scale_1/scale_rename_req
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_scale_1/$exit
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_scale_1/$entry
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_resize_1/index_resize_ack
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_resize_1/index_resize_req
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_resize_1/$exit
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_resize_1/$entry
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_computed_1
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_scaled_1
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_resized_1
      -- 
    req_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(283), ack => array_obj_ref_326_index_offset_req_0); -- 
    access_T_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(60) & access_T_CP_0_elements(123) & access_T_CP_0_elements(280);
      gj_access_T_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	30 
    -- CP-element group 284: marked-predecessors 
    -- CP-element group 284: 	286 
    -- CP-element group 284: 	287 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	286 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_update_start
      -- CP-element group 284: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Update/req
      -- CP-element group 284: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Update/$entry
      -- 
    req_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(284), ack => array_obj_ref_326_index_offset_req_1); -- 
    access_T_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(286) & access_T_CP_0_elements(287);
      gj_access_T_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	283 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	374 
    -- CP-element group 285: marked-successors 
    -- CP-element group 285: 	56 
    -- CP-element group 285: 	119 
    -- CP-element group 285: 	278 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_sample_complete
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Sample/ack
      -- 
    ack_1118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_326_index_offset_ack_0, ack => access_T_CP_0_elements(285)); -- 
    -- CP-element group 286:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	284 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	281 
    -- CP-element group 286: marked-successors 
    -- CP-element group 286: 	284 
    -- CP-element group 286:  members (8) 
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_offset_calculated
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_root_address_calculated
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_base_plus_offset/sum_rename_ack
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_base_plus_offset/sum_rename_req
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_base_plus_offset/$exit
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_base_plus_offset/$entry
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Update/ack
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Update/$exit
      -- 
    ack_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_326_index_offset_ack_1, ack => access_T_CP_0_elements(286)); -- 
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	281 
    -- CP-element group 287: successors 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	281 
    -- CP-element group 287: 	284 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_request/ack
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_request/$exit
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_sample_completed_
      -- 
    ack_1133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_327_final_reg_ack_0, ack => access_T_CP_0_elements(287)); -- 
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	282 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	293 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	282 
    -- CP-element group 288:  members (19) 
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_complete/ack
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_complete/$exit
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_word_addrgen/root_register_req
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_word_addrgen/root_register_ack
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_plus_offset/sum_rename_req
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_word_addrgen/$exit
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_word_addrgen/$entry
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_plus_offset/sum_rename_ack
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_plus_offset/$exit
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_plus_offset/$entry
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_addr_resize/base_resize_ack
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_addr_resize/base_resize_req
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_addr_resize/$exit
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_addr_resize/$entry
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_address_resized
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_root_address_calculated
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_word_address_calculated
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_address_calculated
      -- 
    ack_1138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_327_final_reg_ack_1, ack => access_T_CP_0_elements(288)); -- 
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	60 
    -- CP-element group 289: 	123 
    -- CP-element group 289: 	216 
    -- CP-element group 289: 	280 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Sample/req
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_sample_start_
      -- 
    req_1146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(289), ack => W_fn2_314_delayed_7_0_329_inst_req_0); -- 
    access_T_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(60) & access_T_CP_0_elements(123) & access_T_CP_0_elements(216) & access_T_CP_0_elements(280) & access_T_CP_0_elements(291);
      gj_access_T_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: 	295 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_update_start_
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Update/req
      -- 
    req_1151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(290), ack => W_fn2_314_delayed_7_0_329_inst_req_1); -- 
    access_T_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(292) & access_T_CP_0_elements(295);
      gj_access_T_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	56 
    -- CP-element group 291: 	119 
    -- CP-element group 291: 	212 
    -- CP-element group 291: 	278 
    -- CP-element group 291: 	289 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Sample/$exit
      -- 
    ack_1147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_314_delayed_7_0_329_inst_ack_0, ack => access_T_CP_0_elements(291)); -- 
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	290 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Update/$exit
      -- 
    ack_1152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_314_delayed_7_0_329_inst_ack_1, ack => access_T_CP_0_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	288 
    -- CP-element group 293: 	292 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (5) 
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/word_0/rr
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/word_0/$entry
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/$entry
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/$entry
      -- 
    rr_1185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(293), ack => ptr_deref_335_load_0_req_0); -- 
    access_T_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(288) & access_T_CP_0_elements(292) & access_T_CP_0_elements(295);
      gj_access_T_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	33 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (5) 
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_update_start_
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/word_0/cr
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/word_0/$entry
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/$entry
      -- 
    cr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(294), ack => ptr_deref_335_load_0_req_1); -- 
    access_T_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(296);
      gj_access_T_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	282 
    -- CP-element group 295: 	290 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (5) 
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/word_0/ra
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/word_0/$exit
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/$exit
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/$exit
      -- 
    ra_1186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_335_load_0_ack_0, ack => access_T_CP_0_elements(295)); -- 
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	374 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	154 
    -- CP-element group 296: 	294 
    -- CP-element group 296:  members (9) 
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/word_0/ca
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/word_0/$exit
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/$exit
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/ptr_deref_335_Merge/merge_ack
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/ptr_deref_335_Merge/merge_req
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/ptr_deref_335_Merge/$exit
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/ptr_deref_335_Merge/$entry
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_update_completed_
      -- 
    ca_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_335_load_0_ack_1, ack => access_T_CP_0_elements(296)); -- 
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	60 
    -- CP-element group 297: 	123 
    -- CP-element group 297: 	216 
    -- CP-element group 297: 	280 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Sample/req
      -- CP-element group 297: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_sample_start_
      -- 
    req_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(297), ack => W_fn2_320_delayed_13_0_337_inst_req_0); -- 
    access_T_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(60) & access_T_CP_0_elements(123) & access_T_CP_0_elements(216) & access_T_CP_0_elements(280) & access_T_CP_0_elements(299);
      gj_access_T_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	33 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Update/req
      -- CP-element group 298: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_update_start_
      -- 
    req_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(298), ack => W_fn2_320_delayed_13_0_337_inst_req_1); -- 
    access_T_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(300);
      gj_access_T_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	56 
    -- CP-element group 299: 	119 
    -- CP-element group 299: 	212 
    -- CP-element group 299: 	278 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_sample_completed_
      -- 
    ack_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_320_delayed_13_0_337_inst_ack_0, ack => access_T_CP_0_elements(299)); -- 
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	374 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	154 
    -- CP-element group 300: 	298 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_update_completed_
      -- 
    ack_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_320_delayed_13_0_337_inst_ack_1, ack => access_T_CP_0_elements(300)); -- 
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	159 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Sample/req
      -- CP-element group 301: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Sample/$entry
      -- 
    req_1224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(301), ack => W_fetch_val2_322_delayed_13_0_340_inst_req_0); -- 
    access_T_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(159) & access_T_CP_0_elements(303);
      gj_access_T_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	33 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	304 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Update/req
      -- CP-element group 302: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_update_start_
      -- 
    req_1229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(302), ack => W_fetch_val2_322_delayed_13_0_340_inst_req_1); -- 
    access_T_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(304);
      gj_access_T_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	155 
    -- CP-element group 303: 	301 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_sample_completed_
      -- 
    ack_1225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val2_322_delayed_13_0_340_inst_ack_0, ack => access_T_CP_0_elements(303)); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	374 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	154 
    -- CP-element group 304: 	302 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_update_completed_
      -- 
    ack_1230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val2_322_delayed_13_0_340_inst_ack_1, ack => access_T_CP_0_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	30 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Sample/rr
      -- CP-element group 305: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_sample_start_
      -- 
    rr_1238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(305), ack => type_cast_371_inst_req_0); -- 
    access_T_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(307);
      gj_access_T_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	33 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: 	313 
    -- CP-element group 306: 	319 
    -- CP-element group 306: 	327 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_update_start_
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Update/cr
      -- 
    cr_1243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(306), ack => type_cast_371_inst_req_1); -- 
    access_T_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(308) & access_T_CP_0_elements(313) & access_T_CP_0_elements(319) & access_T_CP_0_elements(327);
      gj_access_T_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Sample/ra
      -- 
    ra_1239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_0, ack => access_T_CP_0_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	311 
    -- CP-element group 308: 	317 
    -- CP-element group 308: 	325 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	76 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Update/ca
      -- 
    ca_1244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_1, ack => access_T_CP_0_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	314 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	315 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	315 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_request/$entry
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_request/req
      -- 
    req_1284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(309), ack => addr_of_399_final_reg_req_0); -- 
    access_T_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(314) & access_T_CP_0_elements(315);
      gj_access_T_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	30 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	316 
    -- CP-element group 310: 	323 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	316 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_update_start_
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_complete/$entry
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_complete/req
      -- 
    req_1289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(310), ack => addr_of_399_final_reg_req_1); -- 
    access_T_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(316) & access_T_CP_0_elements(323);
      gj_access_T_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	81 
    -- CP-element group 311: 	123 
    -- CP-element group 311: 	308 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	313 
    -- CP-element group 311:  members (13) 
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_resized_1
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_scaled_1
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_computed_1
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_resize_1/$entry
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_resize_1/$exit
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_resize_1/index_resize_req
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_resize_1/index_resize_ack
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_scale_1/$entry
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_scale_1/$exit
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_scale_1/scale_rename_req
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_scale_1/scale_rename_ack
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Sample/req
      -- 
    req_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(311), ack => array_obj_ref_398_index_offset_req_0); -- 
    access_T_cp_element_group_311: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_311"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(81) & access_T_CP_0_elements(123) & access_T_CP_0_elements(308);
      gj_access_T_cp_element_group_311 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(311), clk => clk, reset => reset); --
    end block;
    -- CP-element group 312:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	30 
    -- CP-element group 312: marked-predecessors 
    -- CP-element group 312: 	314 
    -- CP-element group 312: 	315 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	314 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_update_start
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Update/req
      -- 
    req_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(312), ack => array_obj_ref_398_index_offset_req_1); -- 
    access_T_cp_element_group_312: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_312"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(314) & access_T_CP_0_elements(315);
      gj_access_T_cp_element_group_312 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(312), clk => clk, reset => reset); --
    end block;
    -- CP-element group 313:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	311 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	374 
    -- CP-element group 313: marked-successors 
    -- CP-element group 313: 	77 
    -- CP-element group 313: 	119 
    -- CP-element group 313: 	306 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_sample_complete
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Sample/ack
      -- 
    ack_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_398_index_offset_ack_0, ack => access_T_CP_0_elements(313)); -- 
    -- CP-element group 314:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	312 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	309 
    -- CP-element group 314: marked-successors 
    -- CP-element group 314: 	312 
    -- CP-element group 314:  members (8) 
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_root_address_calculated
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_offset_calculated
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Update/ack
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_base_plus_offset/$entry
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_base_plus_offset/$exit
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_base_plus_offset/sum_rename_req
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_base_plus_offset/sum_rename_ack
      -- 
    ack_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_398_index_offset_ack_1, ack => access_T_CP_0_elements(314)); -- 
    -- CP-element group 315:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	309 
    -- CP-element group 315: successors 
    -- CP-element group 315: marked-successors 
    -- CP-element group 315: 	309 
    -- CP-element group 315: 	312 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_request/$exit
      -- CP-element group 315: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_request/ack
      -- 
    ack_1285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_399_final_reg_ack_0, ack => access_T_CP_0_elements(315)); -- 
    -- CP-element group 316:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	310 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	321 
    -- CP-element group 316: marked-successors 
    -- CP-element group 316: 	310 
    -- CP-element group 316:  members (19) 
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_complete/$exit
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_complete/ack
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_address_calculated
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_word_address_calculated
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_root_address_calculated
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_address_resized
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_addr_resize/$entry
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_addr_resize/$exit
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_addr_resize/base_resize_req
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_addr_resize/base_resize_ack
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_plus_offset/$entry
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_plus_offset/$exit
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_plus_offset/sum_rename_req
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_plus_offset/sum_rename_ack
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_word_addrgen/$entry
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_word_addrgen/$exit
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_word_addrgen/root_register_req
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_word_addrgen/root_register_ack
      -- 
    ack_1290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_399_final_reg_ack_1, ack => access_T_CP_0_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	81 
    -- CP-element group 317: 	123 
    -- CP-element group 317: 	216 
    -- CP-element group 317: 	308 
    -- CP-element group 317: marked-predecessors 
    -- CP-element group 317: 	319 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	319 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Sample/req
      -- 
    req_1298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(317), ack => W_fn3_374_delayed_7_0_401_inst_req_0); -- 
    access_T_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(81) & access_T_CP_0_elements(123) & access_T_CP_0_elements(216) & access_T_CP_0_elements(308) & access_T_CP_0_elements(319);
      gj_access_T_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: marked-predecessors 
    -- CP-element group 318: 	320 
    -- CP-element group 318: 	323 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	320 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_update_start_
      -- CP-element group 318: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Update/req
      -- 
    req_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(318), ack => W_fn3_374_delayed_7_0_401_inst_req_1); -- 
    access_T_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(320) & access_T_CP_0_elements(323);
      gj_access_T_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	317 
    -- CP-element group 319: successors 
    -- CP-element group 319: marked-successors 
    -- CP-element group 319: 	77 
    -- CP-element group 319: 	119 
    -- CP-element group 319: 	212 
    -- CP-element group 319: 	306 
    -- CP-element group 319: 	317 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Sample/ack
      -- 
    ack_1299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_374_delayed_7_0_401_inst_ack_0, ack => access_T_CP_0_elements(319)); -- 
    -- CP-element group 320:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320: marked-successors 
    -- CP-element group 320: 	318 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_update_completed_
      -- CP-element group 320: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Update/ack
      -- 
    ack_1304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_374_delayed_7_0_401_inst_ack_1, ack => access_T_CP_0_elements(320)); -- 
    -- CP-element group 321:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	316 
    -- CP-element group 321: 	320 
    -- CP-element group 321: marked-predecessors 
    -- CP-element group 321: 	323 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	323 
    -- CP-element group 321:  members (5) 
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_sample_start_
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/$entry
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/$entry
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/word_0/$entry
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/word_0/rr
      -- 
    rr_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(321), ack => ptr_deref_407_load_0_req_0); -- 
    access_T_cp_element_group_321: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_321"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(316) & access_T_CP_0_elements(320) & access_T_CP_0_elements(323);
      gj_access_T_cp_element_group_321 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(321), clk => clk, reset => reset); --
    end block;
    -- CP-element group 322:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	33 
    -- CP-element group 322: marked-predecessors 
    -- CP-element group 322: 	324 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (5) 
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_update_start_
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/$entry
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/$entry
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/word_0/$entry
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/word_0/cr
      -- 
    cr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(322), ack => ptr_deref_407_load_0_req_1); -- 
    access_T_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(324);
      gj_access_T_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: successors 
    -- CP-element group 323: marked-successors 
    -- CP-element group 323: 	310 
    -- CP-element group 323: 	318 
    -- CP-element group 323: 	321 
    -- CP-element group 323:  members (5) 
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/$exit
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/word_0/$exit
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/word_0/ra
      -- 
    ra_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_407_load_0_ack_0, ack => access_T_CP_0_elements(323)); -- 
    -- CP-element group 324:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	374 
    -- CP-element group 324: marked-successors 
    -- CP-element group 324: 	173 
    -- CP-element group 324: 	322 
    -- CP-element group 324:  members (9) 
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/$exit
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/word_0/$exit
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/word_0/ca
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/ptr_deref_407_Merge/$entry
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/ptr_deref_407_Merge/$exit
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/ptr_deref_407_Merge/merge_req
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/ptr_deref_407_Merge/merge_ack
      -- 
    ca_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_407_load_0_ack_1, ack => access_T_CP_0_elements(324)); -- 
    -- CP-element group 325:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	81 
    -- CP-element group 325: 	123 
    -- CP-element group 325: 	216 
    -- CP-element group 325: 	308 
    -- CP-element group 325: marked-predecessors 
    -- CP-element group 325: 	327 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_sample_start_
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Sample/req
      -- 
    req_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(325), ack => W_fn3_380_delayed_13_0_409_inst_req_0); -- 
    access_T_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(81) & access_T_CP_0_elements(123) & access_T_CP_0_elements(216) & access_T_CP_0_elements(308) & access_T_CP_0_elements(327);
      gj_access_T_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	33 
    -- CP-element group 326: marked-predecessors 
    -- CP-element group 326: 	328 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_update_start_
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Update/req
      -- 
    req_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(326), ack => W_fn3_380_delayed_13_0_409_inst_req_1); -- 
    access_T_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(328);
      gj_access_T_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: successors 
    -- CP-element group 327: marked-successors 
    -- CP-element group 327: 	77 
    -- CP-element group 327: 	119 
    -- CP-element group 327: 	212 
    -- CP-element group 327: 	306 
    -- CP-element group 327: 	325 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Sample/ack
      -- 
    ack_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_380_delayed_13_0_409_inst_ack_0, ack => access_T_CP_0_elements(327)); -- 
    -- CP-element group 328:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	374 
    -- CP-element group 328: marked-successors 
    -- CP-element group 328: 	173 
    -- CP-element group 328: 	326 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Update/ack
      -- 
    ack_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_380_delayed_13_0_409_inst_ack_1, ack => access_T_CP_0_elements(328)); -- 
    -- CP-element group 329:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	178 
    -- CP-element group 329: marked-predecessors 
    -- CP-element group 329: 	331 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_sample_start_
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Sample/req
      -- 
    req_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(329), ack => W_fetch_val3_382_delayed_13_0_412_inst_req_0); -- 
    access_T_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(178) & access_T_CP_0_elements(331);
      gj_access_T_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	33 
    -- CP-element group 330: marked-predecessors 
    -- CP-element group 330: 	332 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	332 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_update_start_
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Update/req
      -- 
    req_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(330), ack => W_fetch_val3_382_delayed_13_0_412_inst_req_1); -- 
    access_T_cp_element_group_330: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_330"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(332);
      gj_access_T_cp_element_group_330 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(330), clk => clk, reset => reset); --
    end block;
    -- CP-element group 331:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: successors 
    -- CP-element group 331: marked-successors 
    -- CP-element group 331: 	174 
    -- CP-element group 331: 	329 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Sample/ack
      -- 
    ack_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val3_382_delayed_13_0_412_inst_ack_0, ack => access_T_CP_0_elements(331)); -- 
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	374 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	173 
    -- CP-element group 332: 	330 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Update/ack
      -- 
    ack_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val3_382_delayed_13_0_412_inst_ack_1, ack => access_T_CP_0_elements(332)); -- 
    -- CP-element group 333:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	30 
    -- CP-element group 333: marked-predecessors 
    -- CP-element group 333: 	335 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_sample_start_
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Sample/rr
      -- 
    rr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(333), ack => type_cast_443_inst_req_0); -- 
    access_T_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(335);
      gj_access_T_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	33 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: 	341 
    -- CP-element group 334: 	347 
    -- CP-element group 334: 	355 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_update_start_
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Update/$entry
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Update/cr
      -- 
    cr_1395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(334), ack => type_cast_443_inst_req_1); -- 
    access_T_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(336) & access_T_CP_0_elements(341) & access_T_CP_0_elements(347) & access_T_CP_0_elements(355);
      gj_access_T_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: successors 
    -- CP-element group 335: marked-successors 
    -- CP-element group 335: 	333 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Sample/ra
      -- 
    ra_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_0, ack => access_T_CP_0_elements(335)); -- 
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	339 
    -- CP-element group 336: 	345 
    -- CP-element group 336: 	353 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	97 
    -- CP-element group 336: 	334 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Update/ca
      -- 
    ca_1396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_1, ack => access_T_CP_0_elements(336)); -- 
    -- CP-element group 337:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	342 
    -- CP-element group 337: marked-predecessors 
    -- CP-element group 337: 	343 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	343 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_request/$entry
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_request/req
      -- 
    req_1436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(337), ack => addr_of_471_final_reg_req_0); -- 
    access_T_cp_element_group_337: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_337"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(342) & access_T_CP_0_elements(343);
      gj_access_T_cp_element_group_337 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(337), clk => clk, reset => reset); --
    end block;
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	30 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	344 
    -- CP-element group 338: 	351 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	344 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_update_start_
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_complete/$entry
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_complete/req
      -- 
    req_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(338), ack => addr_of_471_final_reg_req_1); -- 
    access_T_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(344) & access_T_CP_0_elements(351);
      gj_access_T_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	123 
    -- CP-element group 339: 	102 
    -- CP-element group 339: 	336 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (13) 
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_resized_1
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_scaled_1
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_computed_1
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_resize_1/$entry
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_resize_1/$exit
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_resize_1/index_resize_req
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_resize_1/index_resize_ack
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_scale_1/$entry
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_scale_1/$exit
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_scale_1/scale_rename_req
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_scale_1/scale_rename_ack
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Sample/req
      -- 
    req_1421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(339), ack => array_obj_ref_470_index_offset_req_0); -- 
    access_T_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(123) & access_T_CP_0_elements(102) & access_T_CP_0_elements(336);
      gj_access_T_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	30 
    -- CP-element group 340: marked-predecessors 
    -- CP-element group 340: 	342 
    -- CP-element group 340: 	343 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	342 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_update_start
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Update/$entry
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Update/req
      -- 
    req_1426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(340), ack => array_obj_ref_470_index_offset_req_1); -- 
    access_T_cp_element_group_340: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_340"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(342) & access_T_CP_0_elements(343);
      gj_access_T_cp_element_group_340 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(340), clk => clk, reset => reset); --
    end block;
    -- CP-element group 341:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	374 
    -- CP-element group 341: marked-successors 
    -- CP-element group 341: 	119 
    -- CP-element group 341: 	98 
    -- CP-element group 341: 	334 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_sample_complete
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Sample/ack
      -- 
    ack_1422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_470_index_offset_ack_0, ack => access_T_CP_0_elements(341)); -- 
    -- CP-element group 342:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	340 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	337 
    -- CP-element group 342: marked-successors 
    -- CP-element group 342: 	340 
    -- CP-element group 342:  members (8) 
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_root_address_calculated
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_offset_calculated
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_base_plus_offset/$entry
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_base_plus_offset/$exit
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_base_plus_offset/sum_rename_req
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_base_plus_offset/sum_rename_ack
      -- 
    ack_1427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_470_index_offset_ack_1, ack => access_T_CP_0_elements(342)); -- 
    -- CP-element group 343:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	337 
    -- CP-element group 343: successors 
    -- CP-element group 343: marked-successors 
    -- CP-element group 343: 	337 
    -- CP-element group 343: 	340 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_request/$exit
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_request/ack
      -- 
    ack_1437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_471_final_reg_ack_0, ack => access_T_CP_0_elements(343)); -- 
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	338 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	349 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	338 
    -- CP-element group 344:  members (19) 
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_complete/$exit
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_complete/ack
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_address_calculated
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_word_address_calculated
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_root_address_calculated
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_address_resized
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_addr_resize/$entry
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_addr_resize/$exit
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_addr_resize/base_resize_req
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_addr_resize/base_resize_ack
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_plus_offset/$entry
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_plus_offset/$exit
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_plus_offset/sum_rename_req
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_plus_offset/sum_rename_ack
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_word_addrgen/$entry
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_word_addrgen/$exit
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_word_addrgen/root_register_req
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_word_addrgen/root_register_ack
      -- 
    ack_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_471_final_reg_ack_1, ack => access_T_CP_0_elements(344)); -- 
    -- CP-element group 345:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	123 
    -- CP-element group 345: 	102 
    -- CP-element group 345: 	235 
    -- CP-element group 345: 	336 
    -- CP-element group 345: marked-predecessors 
    -- CP-element group 345: 	347 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_sample_start_
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Sample/req
      -- 
    req_1450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(345), ack => W_fn4_434_delayed_7_0_473_inst_req_0); -- 
    access_T_cp_element_group_345: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_345"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(123) & access_T_CP_0_elements(102) & access_T_CP_0_elements(235) & access_T_CP_0_elements(336) & access_T_CP_0_elements(347);
      gj_access_T_cp_element_group_345 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(345), clk => clk, reset => reset); --
    end block;
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	348 
    -- CP-element group 346: 	351 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_update_start_
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Update/$entry
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Update/req
      -- 
    req_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(346), ack => W_fn4_434_delayed_7_0_473_inst_req_1); -- 
    access_T_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(348) & access_T_CP_0_elements(351);
      gj_access_T_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: marked-successors 
    -- CP-element group 347: 	119 
    -- CP-element group 347: 	98 
    -- CP-element group 347: 	231 
    -- CP-element group 347: 	334 
    -- CP-element group 347: 	345 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Sample/ack
      -- 
    ack_1451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn4_434_delayed_7_0_473_inst_ack_0, ack => access_T_CP_0_elements(347)); -- 
    -- CP-element group 348:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348: marked-successors 
    -- CP-element group 348: 	346 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Update/ack
      -- 
    ack_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn4_434_delayed_7_0_473_inst_ack_1, ack => access_T_CP_0_elements(348)); -- 
    -- CP-element group 349:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	344 
    -- CP-element group 349: 	348 
    -- CP-element group 349: marked-predecessors 
    -- CP-element group 349: 	351 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	351 
    -- CP-element group 349:  members (5) 
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_sample_start_
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/$entry
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/word_0/$entry
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/word_0/rr
      -- 
    rr_1489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(349), ack => ptr_deref_479_load_0_req_0); -- 
    access_T_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(344) & access_T_CP_0_elements(348) & access_T_CP_0_elements(351);
      gj_access_T_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	33 
    -- CP-element group 350: marked-predecessors 
    -- CP-element group 350: 	352 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350:  members (5) 
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_update_start_
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/$entry
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/word_0/$entry
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/word_0/cr
      -- 
    cr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(350), ack => ptr_deref_479_load_0_req_1); -- 
    access_T_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(352);
      gj_access_T_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	349 
    -- CP-element group 351: successors 
    -- CP-element group 351: marked-successors 
    -- CP-element group 351: 	338 
    -- CP-element group 351: 	346 
    -- CP-element group 351: 	349 
    -- CP-element group 351:  members (5) 
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_sample_completed_
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/$exit
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/word_0/$exit
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/word_0/ra
      -- 
    ra_1490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_479_load_0_ack_0, ack => access_T_CP_0_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	374 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	192 
    -- CP-element group 352: 	350 
    -- CP-element group 352:  members (9) 
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_update_completed_
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/$exit
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/word_0/$exit
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/word_0/ca
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/ptr_deref_479_Merge/$entry
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/ptr_deref_479_Merge/$exit
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/ptr_deref_479_Merge/merge_req
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/ptr_deref_479_Merge/merge_ack
      -- 
    ca_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_479_load_0_ack_1, ack => access_T_CP_0_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	123 
    -- CP-element group 353: 	102 
    -- CP-element group 353: 	235 
    -- CP-element group 353: 	336 
    -- CP-element group 353: marked-predecessors 
    -- CP-element group 353: 	355 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Sample/req
      -- 
    req_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(353), ack => W_fn4_440_delayed_13_0_481_inst_req_0); -- 
    access_T_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(123) & access_T_CP_0_elements(102) & access_T_CP_0_elements(235) & access_T_CP_0_elements(336) & access_T_CP_0_elements(355);
      gj_access_T_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	33 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_update_start_
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Update/$entry
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Update/req
      -- 
    req_1519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(354), ack => W_fn4_440_delayed_13_0_481_inst_req_1); -- 
    access_T_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(356);
      gj_access_T_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355: marked-successors 
    -- CP-element group 355: 	119 
    -- CP-element group 355: 	98 
    -- CP-element group 355: 	231 
    -- CP-element group 355: 	334 
    -- CP-element group 355: 	353 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Sample/ack
      -- 
    ack_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn4_440_delayed_13_0_481_inst_ack_0, ack => access_T_CP_0_elements(355)); -- 
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	374 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	192 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Update/ack
      -- 
    ack_1520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn4_440_delayed_13_0_481_inst_ack_1, ack => access_T_CP_0_elements(356)); -- 
    -- CP-element group 357:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	197 
    -- CP-element group 357: marked-predecessors 
    -- CP-element group 357: 	359 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_sample_start_
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Sample/$entry
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Sample/req
      -- 
    req_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(357), ack => W_fetch_val4_442_delayed_13_0_484_inst_req_0); -- 
    access_T_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(197) & access_T_CP_0_elements(359);
      gj_access_T_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	33 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_update_start_
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Update/$entry
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Update/req
      -- 
    req_1533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(358), ack => W_fetch_val4_442_delayed_13_0_484_inst_req_1); -- 
    access_T_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(360);
      gj_access_T_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: marked-successors 
    -- CP-element group 359: 	193 
    -- CP-element group 359: 	357 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Sample/ack
      -- 
    ack_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val4_442_delayed_13_0_484_inst_ack_0, ack => access_T_CP_0_elements(359)); -- 
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	374 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	192 
    -- CP-element group 360: 	358 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Update/ack
      -- 
    ack_1534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val4_442_delayed_13_0_484_inst_ack_1, ack => access_T_CP_0_elements(360)); -- 
    -- CP-element group 361:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	140 
    -- CP-element group 361: 	41 
    -- CP-element group 361: 	216 
    -- CP-element group 361: marked-predecessors 
    -- CP-element group 361: 	363 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_sample_start_
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Sample/$entry
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Sample/req
      -- 
    req_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(361), ack => WPIPE_input_pipe1_494_inst_req_0); -- 
    access_T_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(140) & access_T_CP_0_elements(41) & access_T_CP_0_elements(216) & access_T_CP_0_elements(363);
      gj_access_T_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362: marked-successors 
    -- CP-element group 362: 	138 
    -- CP-element group 362: 	37 
    -- CP-element group 362: 	212 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_sample_completed_
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_update_start_
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Sample/ack
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Update/$entry
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Update/req
      -- 
    ack_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_494_inst_ack_0, ack => access_T_CP_0_elements(362)); -- 
    req_1547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(362), ack => WPIPE_input_pipe1_494_inst_req_1); -- 
    -- CP-element group 363:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	374 
    -- CP-element group 363: marked-successors 
    -- CP-element group 363: 	361 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_update_completed_
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Update/ack
      -- 
    ack_1548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_494_inst_ack_1, ack => access_T_CP_0_elements(363)); -- 
    -- CP-element group 364:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	159 
    -- CP-element group 364: 	60 
    -- CP-element group 364: 	216 
    -- CP-element group 364: marked-predecessors 
    -- CP-element group 364: 	366 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_sample_start_
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Sample/$entry
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Sample/req
      -- 
    req_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(364), ack => WPIPE_input_pipe2_498_inst_req_0); -- 
    access_T_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(159) & access_T_CP_0_elements(60) & access_T_CP_0_elements(216) & access_T_CP_0_elements(366);
      gj_access_T_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365: marked-successors 
    -- CP-element group 365: 	155 
    -- CP-element group 365: 	56 
    -- CP-element group 365: 	212 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_update_start_
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Sample/ack
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Update/req
      -- 
    ack_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_498_inst_ack_0, ack => access_T_CP_0_elements(365)); -- 
    req_1561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(365), ack => WPIPE_input_pipe2_498_inst_req_1); -- 
    -- CP-element group 366:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	374 
    -- CP-element group 366: marked-successors 
    -- CP-element group 366: 	364 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Update/ack
      -- 
    ack_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_498_inst_ack_1, ack => access_T_CP_0_elements(366)); -- 
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	81 
    -- CP-element group 367: 	178 
    -- CP-element group 367: 	216 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	369 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_sample_start_
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Sample/$entry
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Sample/req
      -- 
    req_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(367), ack => WPIPE_input_pipe3_502_inst_req_0); -- 
    access_T_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(81) & access_T_CP_0_elements(178) & access_T_CP_0_elements(216) & access_T_CP_0_elements(369);
      gj_access_T_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368: marked-successors 
    -- CP-element group 368: 	77 
    -- CP-element group 368: 	174 
    -- CP-element group 368: 	212 
    -- CP-element group 368:  members (6) 
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_update_start_
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Sample/ack
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Update/req
      -- 
    ack_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_502_inst_ack_0, ack => access_T_CP_0_elements(368)); -- 
    req_1575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(368), ack => WPIPE_input_pipe3_502_inst_req_1); -- 
    -- CP-element group 369:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	374 
    -- CP-element group 369: marked-successors 
    -- CP-element group 369: 	367 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Update/ack
      -- 
    ack_1576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_502_inst_ack_1, ack => access_T_CP_0_elements(369)); -- 
    -- CP-element group 370:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	102 
    -- CP-element group 370: 	197 
    -- CP-element group 370: 	235 
    -- CP-element group 370: marked-predecessors 
    -- CP-element group 370: 	372 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_sample_start_
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Sample/$entry
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Sample/req
      -- 
    req_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(370), ack => WPIPE_input_pipe4_506_inst_req_0); -- 
    access_T_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(102) & access_T_CP_0_elements(197) & access_T_CP_0_elements(235) & access_T_CP_0_elements(372);
      gj_access_T_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371: marked-successors 
    -- CP-element group 371: 	98 
    -- CP-element group 371: 	193 
    -- CP-element group 371: 	231 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_update_start_
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Sample/ack
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Update/$entry
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Update/req
      -- 
    ack_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_506_inst_ack_0, ack => access_T_CP_0_elements(371)); -- 
    req_1589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(371), ack => WPIPE_input_pipe4_506_inst_req_1); -- 
    -- CP-element group 372:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: marked-successors 
    -- CP-element group 372: 	370 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Update/ack
      -- 
    ack_1590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_506_inst_ack_1, ack => access_T_CP_0_elements(372)); -- 
    -- CP-element group 373:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	30 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	31 
    -- CP-element group 373:  members (1) 
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(373) is a control-delay.
    cp_element_373_delay: control_delay_element  generic map(name => " 373_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(30), ack => access_T_CP_0_elements(373), clk => clk, reset =>reset);
    -- CP-element group 374:  join  transition  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	33 
    -- CP-element group 374: 	257 
    -- CP-element group 374: 	268 
    -- CP-element group 374: 	272 
    -- CP-element group 374: 	276 
    -- CP-element group 374: 	285 
    -- CP-element group 374: 	296 
    -- CP-element group 374: 	300 
    -- CP-element group 374: 	304 
    -- CP-element group 374: 	313 
    -- CP-element group 374: 	324 
    -- CP-element group 374: 	328 
    -- CP-element group 374: 	332 
    -- CP-element group 374: 	341 
    -- CP-element group 374: 	352 
    -- CP-element group 374: 	356 
    -- CP-element group 374: 	360 
    -- CP-element group 374: 	363 
    -- CP-element group 374: 	366 
    -- CP-element group 374: 	369 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	27 
    -- CP-element group 374:  members (1) 
      -- CP-element group 374: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/$exit
      -- 
    access_T_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 15,17 => 15,18 => 15,19 => 15,20 => 15);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(257) & access_T_CP_0_elements(268) & access_T_CP_0_elements(272) & access_T_CP_0_elements(276) & access_T_CP_0_elements(285) & access_T_CP_0_elements(296) & access_T_CP_0_elements(300) & access_T_CP_0_elements(304) & access_T_CP_0_elements(313) & access_T_CP_0_elements(324) & access_T_CP_0_elements(328) & access_T_CP_0_elements(332) & access_T_CP_0_elements(341) & access_T_CP_0_elements(352) & access_T_CP_0_elements(356) & access_T_CP_0_elements(360) & access_T_CP_0_elements(363) & access_T_CP_0_elements(366) & access_T_CP_0_elements(369) & access_T_CP_0_elements(372);
      gj_access_T_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  transition  input  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	26 
    -- CP-element group 375: successors 
    -- CP-element group 375:  members (2) 
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_100/loop_exit/$exit
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_100/loop_exit/ack
      -- 
    ack_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_100_branch_ack_0, ack => access_T_CP_0_elements(375)); -- 
    -- CP-element group 376:  transition  input  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	26 
    -- CP-element group 376: successors 
    -- CP-element group 376:  members (2) 
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_100/loop_taken/$exit
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_100/loop_taken/ack
      -- 
    ack_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_100_branch_ack_1, ack => access_T_CP_0_elements(376)); -- 
    -- CP-element group 377:  transition  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	24 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	1 
    -- CP-element group 377:  members (1) 
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_100/$exit
      -- 
    access_T_CP_0_elements(377) <= access_T_CP_0_elements(24);
    access_T_do_while_stmt_100_terminator_1600: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_100_terminator_1600", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(27),loop_continue => access_T_CP_0_elements(376),loop_terminate => access_T_CP_0_elements(375),loop_back => access_T_CP_0_elements(25),loop_exit => access_T_CP_0_elements(24),clk => clk, reset => reset); -- 
    phi_stmt_102_phi_seq_416_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(44);
      access_T_CP_0_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(49);
      access_T_CP_0_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(42);
      access_T_CP_0_elements(51)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(53);
      access_T_CP_0_elements(52)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(54);
      access_T_CP_0_elements(43) <= phi_mux_reqs(1);
      phi_stmt_102_phi_seq_416 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_102_phi_seq_416") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(38), 
          phi_sample_ack => access_T_CP_0_elements(39), 
          phi_update_req => access_T_CP_0_elements(40), 
          phi_update_ack => access_T_CP_0_elements(41), 
          phi_mux_ack => access_T_CP_0_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_107_phi_seq_470_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(63);
      access_T_CP_0_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(70);
      access_T_CP_0_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(71);
      access_T_CP_0_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(61);
      access_T_CP_0_elements(72)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(74);
      access_T_CP_0_elements(73)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(75);
      access_T_CP_0_elements(62) <= phi_mux_reqs(1);
      phi_stmt_107_phi_seq_470 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_107_phi_seq_470") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(57), 
          phi_sample_ack => access_T_CP_0_elements(58), 
          phi_update_req => access_T_CP_0_elements(59), 
          phi_update_ack => access_T_CP_0_elements(60), 
          phi_mux_ack => access_T_CP_0_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_112_phi_seq_524_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(84);
      access_T_CP_0_elements(87)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(91);
      access_T_CP_0_elements(88)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(92);
      access_T_CP_0_elements(85) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(82);
      access_T_CP_0_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(95);
      access_T_CP_0_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(96);
      access_T_CP_0_elements(83) <= phi_mux_reqs(1);
      phi_stmt_112_phi_seq_524 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_112_phi_seq_524") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(78), 
          phi_sample_ack => access_T_CP_0_elements(79), 
          phi_update_req => access_T_CP_0_elements(80), 
          phi_update_ack => access_T_CP_0_elements(81), 
          phi_mux_ack => access_T_CP_0_elements(86), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_117_phi_seq_578_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(105);
      access_T_CP_0_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(112);
      access_T_CP_0_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(113);
      access_T_CP_0_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(103);
      access_T_CP_0_elements(114)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(116);
      access_T_CP_0_elements(115)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(117);
      access_T_CP_0_elements(104) <= phi_mux_reqs(1);
      phi_stmt_117_phi_seq_578 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_117_phi_seq_578") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(99), 
          phi_sample_ack => access_T_CP_0_elements(100), 
          phi_update_req => access_T_CP_0_elements(101), 
          phi_update_ack => access_T_CP_0_elements(102), 
          phi_mux_ack => access_T_CP_0_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_124_phi_seq_622_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(126);
      access_T_CP_0_elements(129)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(129);
      access_T_CP_0_elements(130)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(131);
      access_T_CP_0_elements(127) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(124);
      access_T_CP_0_elements(133)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(134)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(136);
      access_T_CP_0_elements(125) <= phi_mux_reqs(1);
      phi_stmt_124_phi_seq_622 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_124_phi_seq_622") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(120), 
          phi_sample_ack => access_T_CP_0_elements(121), 
          phi_update_req => access_T_CP_0_elements(122), 
          phi_update_ack => access_T_CP_0_elements(123), 
          phi_mux_ack => access_T_CP_0_elements(128), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_129_phi_seq_676_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(143);
      access_T_CP_0_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(148);
      access_T_CP_0_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(149);
      access_T_CP_0_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(141);
      access_T_CP_0_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(152);
      access_T_CP_0_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(153);
      access_T_CP_0_elements(142) <= phi_mux_reqs(1);
      phi_stmt_129_phi_seq_676 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_129_phi_seq_676") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(32), 
          phi_sample_ack => access_T_CP_0_elements(139), 
          phi_update_req => access_T_CP_0_elements(34), 
          phi_update_ack => access_T_CP_0_elements(140), 
          phi_mux_ack => access_T_CP_0_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_133_phi_seq_730_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(162);
      access_T_CP_0_elements(165)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(167);
      access_T_CP_0_elements(166)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(168);
      access_T_CP_0_elements(163) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(160);
      access_T_CP_0_elements(169)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(171);
      access_T_CP_0_elements(170)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(172);
      access_T_CP_0_elements(161) <= phi_mux_reqs(1);
      phi_stmt_133_phi_seq_730 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_133_phi_seq_730") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(156), 
          phi_sample_ack => access_T_CP_0_elements(157), 
          phi_update_req => access_T_CP_0_elements(158), 
          phi_update_ack => access_T_CP_0_elements(159), 
          phi_mux_ack => access_T_CP_0_elements(164), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_137_phi_seq_784_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(181);
      access_T_CP_0_elements(184)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(186);
      access_T_CP_0_elements(185)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(187);
      access_T_CP_0_elements(182) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(179);
      access_T_CP_0_elements(188)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(190);
      access_T_CP_0_elements(189)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(191);
      access_T_CP_0_elements(180) <= phi_mux_reqs(1);
      phi_stmt_137_phi_seq_784 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_137_phi_seq_784") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(175), 
          phi_sample_ack => access_T_CP_0_elements(176), 
          phi_update_req => access_T_CP_0_elements(177), 
          phi_update_ack => access_T_CP_0_elements(178), 
          phi_mux_ack => access_T_CP_0_elements(183), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_141_phi_seq_838_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(200);
      access_T_CP_0_elements(203)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(205);
      access_T_CP_0_elements(204)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(206);
      access_T_CP_0_elements(201) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(198);
      access_T_CP_0_elements(207)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(209);
      access_T_CP_0_elements(208)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(210);
      access_T_CP_0_elements(199) <= phi_mux_reqs(1);
      phi_stmt_141_phi_seq_838 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_141_phi_seq_838") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(194), 
          phi_sample_ack => access_T_CP_0_elements(195), 
          phi_update_req => access_T_CP_0_elements(196), 
          phi_update_ack => access_T_CP_0_elements(197), 
          phi_mux_ack => access_T_CP_0_elements(202), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_145_phi_seq_882_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(219);
      access_T_CP_0_elements(222)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(222);
      access_T_CP_0_elements(223)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(224);
      access_T_CP_0_elements(220) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(217);
      access_T_CP_0_elements(226)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(228);
      access_T_CP_0_elements(227)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(229);
      access_T_CP_0_elements(218) <= phi_mux_reqs(1);
      phi_stmt_145_phi_seq_882 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_145_phi_seq_882") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(213), 
          phi_sample_ack => access_T_CP_0_elements(214), 
          phi_update_req => access_T_CP_0_elements(215), 
          phi_update_ack => access_T_CP_0_elements(216), 
          phi_mux_ack => access_T_CP_0_elements(221), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_150_phi_seq_926_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(238);
      access_T_CP_0_elements(241)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(241);
      access_T_CP_0_elements(242)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(243);
      access_T_CP_0_elements(239) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(236);
      access_T_CP_0_elements(245)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(247);
      access_T_CP_0_elements(246)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(248);
      access_T_CP_0_elements(237) <= phi_mux_reqs(1);
      phi_stmt_150_phi_seq_926 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_150_phi_seq_926") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(232), 
          phi_sample_ack => access_T_CP_0_elements(233), 
          phi_update_req => access_T_CP_0_elements(234), 
          phi_update_ack => access_T_CP_0_elements(235), 
          phi_mux_ack => access_T_CP_0_elements(240), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_368_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(28);
        preds(1)  <= access_T_CP_0_elements(29);
        entry_tmerge_368 : transition_merge -- 
          generic map(name => " entry_tmerge_368")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(30));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_183_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_191_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_121_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_166_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_91_wire : std_logic_vector(31 downto 0);
    signal ADD_u64_u64_233_wire : std_logic_vector(63 downto 0);
    signal ADD_u64_u64_305_wire : std_logic_vector(63 downto 0);
    signal ADD_u64_u64_377_wire : std_logic_vector(63 downto 0);
    signal ADD_u64_u64_449_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_209_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_281_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_353_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_425_wire : std_logic_vector(63 downto 0);
    signal LSHR_u32_u32_59_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_73_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_87_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_90_wire : std_logic_vector(31 downto 0);
    signal LSHR_u64_u64_217_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_240_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_243_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_253_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_253_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_253_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_289_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_312_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_315_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_325_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_325_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_325_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_361_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_384_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_387_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_397_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_397_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_397_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_433_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_456_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_459_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_469_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_469_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_469_wire : std_logic_vector(63 downto 0);
    signal MUL_u16_u16_34_wire : std_logic_vector(15 downto 0);
    signal NEQ_u64_u1_244_wire : std_logic_vector(0 downto 0);
    signal NEQ_u64_u1_316_wire : std_logic_vector(0 downto 0);
    signal NEQ_u64_u1_388_wire : std_logic_vector(0 downto 0);
    signal NEQ_u64_u1_460_wire : std_logic_vector(0 downto 0);
    signal SUB_u64_u64_210_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_282_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_354_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_426_wire : std_logic_vector(63 downto 0);
    signal address1_102 : std_logic_vector(63 downto 0);
    signal address2_107 : std_logic_vector(63 downto 0);
    signal address3_112 : std_logic_vector(63 downto 0);
    signal address4_117 : std_logic_vector(63 downto 0);
    signal array_obj_ref_254_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_254_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_254_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_254_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_254_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_254_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_root_address : std_logic_vector(13 downto 0);
    signal continue1_199 : std_logic_vector(0 downto 0);
    signal continue2_204 : std_logic_vector(0 downto 0);
    signal fetch_add1_49 : std_logic_vector(31 downto 0);
    signal fetch_add2_63 : std_logic_vector(31 downto 0);
    signal fetch_add3_77 : std_logic_vector(31 downto 0);
    signal fetch_add4_95 : std_logic_vector(31 downto 0);
    signal fetch_addr1_256 : std_logic_vector(31 downto 0);
    signal fetch_addr2_328 : std_logic_vector(31 downto 0);
    signal fetch_addr3_400 : std_logic_vector(31 downto 0);
    signal fetch_addr4_472 : std_logic_vector(31 downto 0);
    signal fetch_val1_129 : std_logic_vector(63 downto 0);
    signal fetch_val1_262_delayed_13_0_270 : std_logic_vector(63 downto 0);
    signal fetch_val2_133 : std_logic_vector(63 downto 0);
    signal fetch_val2_322_delayed_13_0_342 : std_logic_vector(63 downto 0);
    signal fetch_val3_137 : std_logic_vector(63 downto 0);
    signal fetch_val3_382_delayed_13_0_414 : std_logic_vector(63 downto 0);
    signal fetch_val4_141 : std_logic_vector(63 downto 0);
    signal fetch_val4_442_delayed_13_0_486 : std_logic_vector(63 downto 0);
    signal fn1_247 : std_logic_vector(0 downto 0);
    signal fn1_254_delayed_7_0_259 : std_logic_vector(0 downto 0);
    signal fn1_260_delayed_13_0_267 : std_logic_vector(0 downto 0);
    signal fn2_314_delayed_7_0_331 : std_logic_vector(0 downto 0);
    signal fn2_319 : std_logic_vector(0 downto 0);
    signal fn2_320_delayed_13_0_339 : std_logic_vector(0 downto 0);
    signal fn3_374_delayed_7_0_403 : std_logic_vector(0 downto 0);
    signal fn3_380_delayed_13_0_411 : std_logic_vector(0 downto 0);
    signal fn3_391 : std_logic_vector(0 downto 0);
    signal fn4_434_delayed_7_0_475 : std_logic_vector(0 downto 0);
    signal fn4_440_delayed_13_0_483 : std_logic_vector(0 downto 0);
    signal fn4_463 : std_logic_vector(0 downto 0);
    signal fv1_264 : std_logic_vector(63 downto 0);
    signal fv2_336 : std_logic_vector(63 downto 0);
    signal fv3_408 : std_logic_vector(63 downto 0);
    signal fv4_480 : std_logic_vector(63 downto 0);
    signal konst_163_wire_constant : std_logic_vector(31 downto 0);
    signal konst_165_wire_constant : std_logic_vector(31 downto 0);
    signal konst_182_wire_constant : std_logic_vector(15 downto 0);
    signal konst_190_wire_constant : std_logic_vector(15 downto 0);
    signal konst_206_wire_constant : std_logic_vector(63 downto 0);
    signal konst_208_wire_constant : std_logic_vector(63 downto 0);
    signal konst_211_wire_constant : std_logic_vector(63 downto 0);
    signal konst_222_wire_constant : std_logic_vector(63 downto 0);
    signal konst_239_wire_constant : std_logic_vector(63 downto 0);
    signal konst_242_wire_constant : std_logic_vector(63 downto 0);
    signal konst_252_wire_constant : std_logic_vector(63 downto 0);
    signal konst_278_wire_constant : std_logic_vector(63 downto 0);
    signal konst_280_wire_constant : std_logic_vector(63 downto 0);
    signal konst_283_wire_constant : std_logic_vector(63 downto 0);
    signal konst_294_wire_constant : std_logic_vector(63 downto 0);
    signal konst_311_wire_constant : std_logic_vector(63 downto 0);
    signal konst_314_wire_constant : std_logic_vector(63 downto 0);
    signal konst_324_wire_constant : std_logic_vector(63 downto 0);
    signal konst_350_wire_constant : std_logic_vector(63 downto 0);
    signal konst_352_wire_constant : std_logic_vector(63 downto 0);
    signal konst_355_wire_constant : std_logic_vector(63 downto 0);
    signal konst_366_wire_constant : std_logic_vector(63 downto 0);
    signal konst_383_wire_constant : std_logic_vector(63 downto 0);
    signal konst_386_wire_constant : std_logic_vector(63 downto 0);
    signal konst_396_wire_constant : std_logic_vector(63 downto 0);
    signal konst_39_wire_constant : std_logic_vector(31 downto 0);
    signal konst_422_wire_constant : std_logic_vector(63 downto 0);
    signal konst_424_wire_constant : std_logic_vector(63 downto 0);
    signal konst_427_wire_constant : std_logic_vector(63 downto 0);
    signal konst_438_wire_constant : std_logic_vector(63 downto 0);
    signal konst_455_wire_constant : std_logic_vector(63 downto 0);
    signal konst_458_wire_constant : std_logic_vector(63 downto 0);
    signal konst_468_wire_constant : std_logic_vector(63 downto 0);
    signal konst_58_wire_constant : std_logic_vector(31 downto 0);
    signal konst_72_wire_constant : std_logic_vector(31 downto 0);
    signal konst_86_wire_constant : std_logic_vector(31 downto 0);
    signal konst_89_wire_constant : std_logic_vector(31 downto 0);
    signal m2_factor_41 : std_logic_vector(31 downto 0);
    signal m_factor_36 : std_logic_vector(31 downto 0);
    signal my_fetch1_53 : std_logic_vector(63 downto 0);
    signal my_fetch1_53_131_buffered : std_logic_vector(63 downto 0);
    signal my_fetch2_67 : std_logic_vector(63 downto 0);
    signal my_fetch2_67_135_buffered : std_logic_vector(63 downto 0);
    signal my_fetch3_81 : std_logic_vector(63 downto 0);
    signal my_fetch3_81_139_buffered : std_logic_vector(63 downto 0);
    signal my_fetch4_99 : std_logic_vector(63 downto 0);
    signal my_fetch4_99_143_buffered : std_logic_vector(63 downto 0);
    signal my_num1_213 : std_logic_vector(63 downto 0);
    signal my_num2_285 : std_logic_vector(63 downto 0);
    signal my_num3_357 : std_logic_vector(63 downto 0);
    signal my_num4_429 : std_logic_vector(63 downto 0);
    signal mycounter_124 : std_logic_vector(31 downto 0);
    signal n_address1_236 : std_logic_vector(63 downto 0);
    signal n_address1_236_106_buffered : std_logic_vector(63 downto 0);
    signal n_address2_308 : std_logic_vector(63 downto 0);
    signal n_address2_308_111_buffered : std_logic_vector(63 downto 0);
    signal n_address3_380 : std_logic_vector(63 downto 0);
    signal n_address3_380_116_buffered : std_logic_vector(63 downto 0);
    signal n_address4_452 : std_logic_vector(63 downto 0);
    signal n_address4_452_123_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val1_276 : std_logic_vector(63 downto 0);
    signal n_fetch_val1_276_132_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val2_348 : std_logic_vector(63 downto 0);
    signal n_fetch_val2_348_136_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val3_420 : std_logic_vector(63 downto 0);
    signal n_fetch_val3_420_140_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val4_492 : std_logic_vector(63 downto 0);
    signal n_fetch_val4_492_144_buffered : std_logic_vector(63 downto 0);
    signal n_mycounter_168 : std_logic_vector(31 downto 0);
    signal n_mycounter_168_128_buffered : std_logic_vector(31 downto 0);
    signal n_row1_186 : std_logic_vector(15 downto 0);
    signal n_row1_186_149_buffered : std_logic_vector(15 downto 0);
    signal n_row2_194 : std_logic_vector(15 downto 0);
    signal n_row2_194_154_buffered : std_logic_vector(15 downto 0);
    signal next_row_160 : std_logic_vector(0 downto 0);
    signal ptr_deref_263_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_263_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_263_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_263_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_263_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_335_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_335_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_335_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_335_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_335_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_407_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_407_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_407_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_407_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_407_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_479_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_479_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_479_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_479_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_479_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_52_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_52_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_52_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_52_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_52_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_66_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_66_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_66_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_66_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_66_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_80_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_80_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_80_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_80_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_80_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_98_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_98_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_98_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_98_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_98_word_offset_0 : std_logic_vector(13 downto 0);
    signal row1_145 : std_logic_vector(15 downto 0);
    signal row2_150 : std_logic_vector(15 downto 0);
    signal send_now1_173 : std_logic_vector(0 downto 0);
    signal send_now2_178 : std_logic_vector(0 downto 0);
    signal temp_address1_224 : std_logic_vector(63 downto 0);
    signal temp_address2_296 : std_logic_vector(63 downto 0);
    signal temp_address3_368 : std_logic_vector(63 downto 0);
    signal temp_address4_440 : std_logic_vector(63 downto 0);
    signal type_cast_105_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_110_wire : std_logic_vector(63 downto 0);
    signal type_cast_115_wire : std_logic_vector(63 downto 0);
    signal type_cast_122_wire : std_logic_vector(63 downto 0);
    signal type_cast_127_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_148_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_153_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_229_229_delayed_1_0_228 : std_logic_vector(63 downto 0);
    signal type_cast_289_289_delayed_1_0_300 : std_logic_vector(63 downto 0);
    signal type_cast_349_349_delayed_1_0_372 : std_logic_vector(63 downto 0);
    signal type_cast_409_409_delayed_1_0_444 : std_logic_vector(63 downto 0);
    signal type_cast_60_resized : std_logic_vector(13 downto 0);
    signal type_cast_60_scaled : std_logic_vector(13 downto 0);
    signal type_cast_60_wire : std_logic_vector(63 downto 0);
    signal type_cast_74_resized : std_logic_vector(13 downto 0);
    signal type_cast_74_scaled : std_logic_vector(13 downto 0);
    signal type_cast_74_wire : std_logic_vector(63 downto 0);
    signal type_cast_92_resized : std_logic_vector(13 downto 0);
    signal type_cast_92_scaled : std_logic_vector(13 downto 0);
    signal type_cast_92_wire : std_logic_vector(63 downto 0);
    signal var_val1_219 : std_logic_vector(7 downto 0);
    signal var_val2_291 : std_logic_vector(7 downto 0);
    signal var_val3_363 : std_logic_vector(7 downto 0);
    signal var_val4_435 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_254_constant_part_of_offset <= "00000000000000";
    array_obj_ref_254_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_254_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_254_resized_base_address <= "00000000000000";
    array_obj_ref_326_constant_part_of_offset <= "00000000000000";
    array_obj_ref_326_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_326_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_326_resized_base_address <= "00000000000000";
    array_obj_ref_398_constant_part_of_offset <= "00000000000000";
    array_obj_ref_398_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_398_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_398_resized_base_address <= "00000000000000";
    array_obj_ref_470_constant_part_of_offset <= "00000000000000";
    array_obj_ref_470_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_470_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_470_resized_base_address <= "00000000000000";
    array_obj_ref_61_constant_part_of_offset <= "00000000000000";
    array_obj_ref_61_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_61_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_61_resized_base_address <= "00000000000000";
    array_obj_ref_75_constant_part_of_offset <= "00000000000000";
    array_obj_ref_75_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_75_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_75_resized_base_address <= "00000000000000";
    array_obj_ref_93_constant_part_of_offset <= "00000000000000";
    array_obj_ref_93_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_93_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_93_resized_base_address <= "00000000000000";
    fetch_add1_49 <= "00000000000000000000000000000000";
    konst_163_wire_constant <= "00000000000000000000000000000001";
    konst_165_wire_constant <= "00000000000000000000000000000001";
    konst_182_wire_constant <= "0000000000000010";
    konst_190_wire_constant <= "0000000000000010";
    konst_206_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_208_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_211_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_222_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_239_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_242_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_252_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_278_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_280_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_283_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_294_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_311_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_314_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_324_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_350_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_352_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_355_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_366_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_383_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_396_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_39_wire_constant <= "00000000000000000000000000000001";
    konst_422_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_424_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_427_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_438_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_455_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_458_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_468_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_58_wire_constant <= "00000000000000000000000000000011";
    konst_72_wire_constant <= "00000000000000000000000000000010";
    konst_86_wire_constant <= "00000000000000000000000000000010";
    konst_89_wire_constant <= "00000000000000000000000000000011";
    ptr_deref_263_word_offset_0 <= "00000000000000";
    ptr_deref_335_word_offset_0 <= "00000000000000";
    ptr_deref_407_word_offset_0 <= "00000000000000";
    ptr_deref_479_word_offset_0 <= "00000000000000";
    ptr_deref_52_word_offset_0 <= "00000000000000";
    ptr_deref_66_word_offset_0 <= "00000000000000";
    ptr_deref_80_word_offset_0 <= "00000000000000";
    ptr_deref_98_word_offset_0 <= "00000000000000";
    type_cast_105_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_127_wire_constant <= "00000000000000000000000000000001";
    type_cast_148_wire_constant <= "0000000000000000";
    type_cast_153_wire_constant <= "0000000000000001";
    phi_stmt_102: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_105_wire_constant & n_address1_236_106_buffered;
      req <= phi_stmt_102_req_0 & phi_stmt_102_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_102",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_102_ack_0,
          idata => idata,
          odata => address1_102,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_102
    phi_stmt_107: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_110_wire & n_address2_308_111_buffered;
      req <= phi_stmt_107_req_0 & phi_stmt_107_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_107",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_107_ack_0,
          idata => idata,
          odata => address2_107,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_107
    phi_stmt_112: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_115_wire & n_address3_380_116_buffered;
      req <= phi_stmt_112_req_0 & phi_stmt_112_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_112",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_112_ack_0,
          idata => idata,
          odata => address3_112,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_112
    phi_stmt_117: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_122_wire & n_address4_452_123_buffered;
      req <= phi_stmt_117_req_0 & phi_stmt_117_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_117",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_117_ack_0,
          idata => idata,
          odata => address4_117,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_117
    phi_stmt_124: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_127_wire_constant & n_mycounter_168_128_buffered;
      req <= phi_stmt_124_req_0 & phi_stmt_124_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_124",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_124_ack_0,
          idata => idata,
          odata => mycounter_124,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_124
    phi_stmt_129: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch1_53_131_buffered & n_fetch_val1_276_132_buffered;
      req <= phi_stmt_129_req_0 & phi_stmt_129_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_129",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_129_ack_0,
          idata => idata,
          odata => fetch_val1_129,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_129
    phi_stmt_133: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch2_67_135_buffered & n_fetch_val2_348_136_buffered;
      req <= phi_stmt_133_req_0 & phi_stmt_133_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_133",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_133_ack_0,
          idata => idata,
          odata => fetch_val2_133,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_133
    phi_stmt_137: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch3_81_139_buffered & n_fetch_val3_420_140_buffered;
      req <= phi_stmt_137_req_0 & phi_stmt_137_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_137",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_137_ack_0,
          idata => idata,
          odata => fetch_val3_137,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_137
    phi_stmt_141: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch4_99_143_buffered & n_fetch_val4_492_144_buffered;
      req <= phi_stmt_141_req_0 & phi_stmt_141_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_141",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_141_ack_0,
          idata => idata,
          odata => fetch_val4_141,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_141
    phi_stmt_145: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_148_wire_constant & n_row1_186_149_buffered;
      req <= phi_stmt_145_req_0 & phi_stmt_145_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_145",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_145_ack_0,
          idata => idata,
          odata => row1_145,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_145
    phi_stmt_150: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_153_wire_constant & n_row2_194_154_buffered;
      req <= phi_stmt_150_req_0 & phi_stmt_150_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_150",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_150_ack_0,
          idata => idata,
          odata => row2_150,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_150
    -- flow-through select operator MUX_167_inst
    n_mycounter_168 <= konst_163_wire_constant when (next_row_160(0) /=  '0') else ADD_u32_u32_166_wire;
    -- flow-through select operator MUX_185_inst
    n_row1_186 <= ADD_u16_u16_183_wire when (next_row_160(0) /=  '0') else row1_145;
    -- flow-through select operator MUX_193_inst
    n_row2_194 <= ADD_u16_u16_191_wire when (next_row_160(0) /=  '0') else row2_150;
    -- flow-through select operator MUX_235_inst
    n_address1_236 <= ADD_u64_u64_233_wire when (next_row_160(0) /=  '0') else temp_address1_224;
    -- flow-through select operator MUX_275_inst
    n_fetch_val1_276 <= fv1_264 when (fn1_260_delayed_13_0_267(0) /=  '0') else fetch_val1_262_delayed_13_0_270;
    -- flow-through select operator MUX_307_inst
    n_address2_308 <= ADD_u64_u64_305_wire when (next_row_160(0) /=  '0') else temp_address2_296;
    -- flow-through select operator MUX_347_inst
    n_fetch_val2_348 <= fv2_336 when (fn2_320_delayed_13_0_339(0) /=  '0') else fetch_val2_322_delayed_13_0_342;
    -- flow-through select operator MUX_379_inst
    n_address3_380 <= ADD_u64_u64_377_wire when (next_row_160(0) /=  '0') else temp_address3_368;
    -- flow-through select operator MUX_419_inst
    n_fetch_val3_420 <= fv3_408 when (fn3_380_delayed_13_0_411(0) /=  '0') else fetch_val3_382_delayed_13_0_414;
    -- flow-through select operator MUX_451_inst
    n_address4_452 <= ADD_u64_u64_449_wire when (next_row_160(0) /=  '0') else temp_address4_440;
    -- flow-through select operator MUX_491_inst
    n_fetch_val4_492 <= fv4_480 when (fn4_440_delayed_13_0_483(0) /=  '0') else fetch_val4_442_delayed_13_0_486;
    W_fetch_val1_262_delayed_13_0_268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val1_262_delayed_13_0_268_inst_req_0;
      W_fetch_val1_262_delayed_13_0_268_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val1_262_delayed_13_0_268_inst_req_1;
      W_fetch_val1_262_delayed_13_0_268_inst_ack_1<= rack(0);
      W_fetch_val1_262_delayed_13_0_268_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val1_262_delayed_13_0_268_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val1_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val1_262_delayed_13_0_270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val2_322_delayed_13_0_340_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val2_322_delayed_13_0_340_inst_req_0;
      W_fetch_val2_322_delayed_13_0_340_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val2_322_delayed_13_0_340_inst_req_1;
      W_fetch_val2_322_delayed_13_0_340_inst_ack_1<= rack(0);
      W_fetch_val2_322_delayed_13_0_340_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val2_322_delayed_13_0_340_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val2_133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val2_322_delayed_13_0_342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val3_382_delayed_13_0_412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val3_382_delayed_13_0_412_inst_req_0;
      W_fetch_val3_382_delayed_13_0_412_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val3_382_delayed_13_0_412_inst_req_1;
      W_fetch_val3_382_delayed_13_0_412_inst_ack_1<= rack(0);
      W_fetch_val3_382_delayed_13_0_412_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val3_382_delayed_13_0_412_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val3_137,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val3_382_delayed_13_0_414,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val4_442_delayed_13_0_484_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val4_442_delayed_13_0_484_inst_req_0;
      W_fetch_val4_442_delayed_13_0_484_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val4_442_delayed_13_0_484_inst_req_1;
      W_fetch_val4_442_delayed_13_0_484_inst_ack_1<= rack(0);
      W_fetch_val4_442_delayed_13_0_484_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val4_442_delayed_13_0_484_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val4_141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val4_442_delayed_13_0_486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn1_254_delayed_7_0_257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn1_254_delayed_7_0_257_inst_req_0;
      W_fn1_254_delayed_7_0_257_inst_ack_0<= wack(0);
      rreq(0) <= W_fn1_254_delayed_7_0_257_inst_req_1;
      W_fn1_254_delayed_7_0_257_inst_ack_1<= rack(0);
      W_fn1_254_delayed_7_0_257_inst : InterlockBuffer generic map ( -- 
        name => "W_fn1_254_delayed_7_0_257_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn1_247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn1_254_delayed_7_0_259,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn1_260_delayed_13_0_265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn1_260_delayed_13_0_265_inst_req_0;
      W_fn1_260_delayed_13_0_265_inst_ack_0<= wack(0);
      rreq(0) <= W_fn1_260_delayed_13_0_265_inst_req_1;
      W_fn1_260_delayed_13_0_265_inst_ack_1<= rack(0);
      W_fn1_260_delayed_13_0_265_inst : InterlockBuffer generic map ( -- 
        name => "W_fn1_260_delayed_13_0_265_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn1_247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn1_260_delayed_13_0_267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn2_314_delayed_7_0_329_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn2_314_delayed_7_0_329_inst_req_0;
      W_fn2_314_delayed_7_0_329_inst_ack_0<= wack(0);
      rreq(0) <= W_fn2_314_delayed_7_0_329_inst_req_1;
      W_fn2_314_delayed_7_0_329_inst_ack_1<= rack(0);
      W_fn2_314_delayed_7_0_329_inst : InterlockBuffer generic map ( -- 
        name => "W_fn2_314_delayed_7_0_329_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn2_319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn2_314_delayed_7_0_331,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn2_320_delayed_13_0_337_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn2_320_delayed_13_0_337_inst_req_0;
      W_fn2_320_delayed_13_0_337_inst_ack_0<= wack(0);
      rreq(0) <= W_fn2_320_delayed_13_0_337_inst_req_1;
      W_fn2_320_delayed_13_0_337_inst_ack_1<= rack(0);
      W_fn2_320_delayed_13_0_337_inst : InterlockBuffer generic map ( -- 
        name => "W_fn2_320_delayed_13_0_337_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn2_319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn2_320_delayed_13_0_339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn3_374_delayed_7_0_401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn3_374_delayed_7_0_401_inst_req_0;
      W_fn3_374_delayed_7_0_401_inst_ack_0<= wack(0);
      rreq(0) <= W_fn3_374_delayed_7_0_401_inst_req_1;
      W_fn3_374_delayed_7_0_401_inst_ack_1<= rack(0);
      W_fn3_374_delayed_7_0_401_inst : InterlockBuffer generic map ( -- 
        name => "W_fn3_374_delayed_7_0_401_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn3_391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn3_374_delayed_7_0_403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn3_380_delayed_13_0_409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn3_380_delayed_13_0_409_inst_req_0;
      W_fn3_380_delayed_13_0_409_inst_ack_0<= wack(0);
      rreq(0) <= W_fn3_380_delayed_13_0_409_inst_req_1;
      W_fn3_380_delayed_13_0_409_inst_ack_1<= rack(0);
      W_fn3_380_delayed_13_0_409_inst : InterlockBuffer generic map ( -- 
        name => "W_fn3_380_delayed_13_0_409_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn3_391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn3_380_delayed_13_0_411,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn4_434_delayed_7_0_473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn4_434_delayed_7_0_473_inst_req_0;
      W_fn4_434_delayed_7_0_473_inst_ack_0<= wack(0);
      rreq(0) <= W_fn4_434_delayed_7_0_473_inst_req_1;
      W_fn4_434_delayed_7_0_473_inst_ack_1<= rack(0);
      W_fn4_434_delayed_7_0_473_inst : InterlockBuffer generic map ( -- 
        name => "W_fn4_434_delayed_7_0_473_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn4_463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn4_434_delayed_7_0_475,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn4_440_delayed_13_0_481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn4_440_delayed_13_0_481_inst_req_0;
      W_fn4_440_delayed_13_0_481_inst_ack_0<= wack(0);
      rreq(0) <= W_fn4_440_delayed_13_0_481_inst_req_1;
      W_fn4_440_delayed_13_0_481_inst_ack_1<= rack(0);
      W_fn4_440_delayed_13_0_481_inst : InterlockBuffer generic map ( -- 
        name => "W_fn4_440_delayed_13_0_481_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn4_463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn4_440_delayed_13_0_483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_255_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_255_final_reg_req_0;
      addr_of_255_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_255_final_reg_req_1;
      addr_of_255_final_reg_ack_1<= rack(0);
      addr_of_255_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_255_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_254_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_327_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_327_final_reg_req_0;
      addr_of_327_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_327_final_reg_req_1;
      addr_of_327_final_reg_ack_1<= rack(0);
      addr_of_327_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_327_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_326_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_328,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_399_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_399_final_reg_req_0;
      addr_of_399_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_399_final_reg_req_1;
      addr_of_399_final_reg_ack_1<= rack(0);
      addr_of_399_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_399_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_398_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr3_400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_471_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_471_final_reg_req_0;
      addr_of_471_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_471_final_reg_req_1;
      addr_of_471_final_reg_ack_1<= rack(0);
      addr_of_471_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_471_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_470_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr4_472,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_62_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_62_final_reg_req_0;
      addr_of_62_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_62_final_reg_req_1;
      addr_of_62_final_reg_ack_1<= rack(0);
      addr_of_62_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_62_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_61_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_add2_63,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_76_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_76_final_reg_req_0;
      addr_of_76_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_76_final_reg_req_1;
      addr_of_76_final_reg_ack_1<= rack(0);
      addr_of_76_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_76_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_75_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_add3_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_94_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_94_final_reg_req_0;
      addr_of_94_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_94_final_reg_req_1;
      addr_of_94_final_reg_ack_1<= rack(0);
      addr_of_94_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_94_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_93_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_add4_95,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch1_53_131_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch1_53_131_buf_req_0;
      my_fetch1_53_131_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch1_53_131_buf_req_1;
      my_fetch1_53_131_buf_ack_1<= rack(0);
      my_fetch1_53_131_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch1_53_131_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch1_53,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch1_53_131_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch2_67_135_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch2_67_135_buf_req_0;
      my_fetch2_67_135_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch2_67_135_buf_req_1;
      my_fetch2_67_135_buf_ack_1<= rack(0);
      my_fetch2_67_135_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch2_67_135_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch2_67,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch2_67_135_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch3_81_139_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch3_81_139_buf_req_0;
      my_fetch3_81_139_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch3_81_139_buf_req_1;
      my_fetch3_81_139_buf_ack_1<= rack(0);
      my_fetch3_81_139_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch3_81_139_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch3_81,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch3_81_139_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch4_99_143_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch4_99_143_buf_req_0;
      my_fetch4_99_143_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch4_99_143_buf_req_1;
      my_fetch4_99_143_buf_ack_1<= rack(0);
      my_fetch4_99_143_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch4_99_143_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch4_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch4_99_143_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address1_236_106_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address1_236_106_buf_req_0;
      n_address1_236_106_buf_ack_0<= wack(0);
      rreq(0) <= n_address1_236_106_buf_req_1;
      n_address1_236_106_buf_ack_1<= rack(0);
      n_address1_236_106_buf : InterlockBuffer generic map ( -- 
        name => "n_address1_236_106_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address1_236,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address1_236_106_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address2_308_111_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address2_308_111_buf_req_0;
      n_address2_308_111_buf_ack_0<= wack(0);
      rreq(0) <= n_address2_308_111_buf_req_1;
      n_address2_308_111_buf_ack_1<= rack(0);
      n_address2_308_111_buf : InterlockBuffer generic map ( -- 
        name => "n_address2_308_111_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address2_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address2_308_111_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address3_380_116_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address3_380_116_buf_req_0;
      n_address3_380_116_buf_ack_0<= wack(0);
      rreq(0) <= n_address3_380_116_buf_req_1;
      n_address3_380_116_buf_ack_1<= rack(0);
      n_address3_380_116_buf : InterlockBuffer generic map ( -- 
        name => "n_address3_380_116_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address3_380,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address3_380_116_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address4_452_123_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address4_452_123_buf_req_0;
      n_address4_452_123_buf_ack_0<= wack(0);
      rreq(0) <= n_address4_452_123_buf_req_1;
      n_address4_452_123_buf_ack_1<= rack(0);
      n_address4_452_123_buf : InterlockBuffer generic map ( -- 
        name => "n_address4_452_123_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address4_452,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address4_452_123_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val1_276_132_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val1_276_132_buf_req_0;
      n_fetch_val1_276_132_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val1_276_132_buf_req_1;
      n_fetch_val1_276_132_buf_ack_1<= rack(0);
      n_fetch_val1_276_132_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val1_276_132_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val1_276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val1_276_132_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val2_348_136_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val2_348_136_buf_req_0;
      n_fetch_val2_348_136_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val2_348_136_buf_req_1;
      n_fetch_val2_348_136_buf_ack_1<= rack(0);
      n_fetch_val2_348_136_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val2_348_136_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val2_348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val2_348_136_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val3_420_140_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val3_420_140_buf_req_0;
      n_fetch_val3_420_140_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val3_420_140_buf_req_1;
      n_fetch_val3_420_140_buf_ack_1<= rack(0);
      n_fetch_val3_420_140_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val3_420_140_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val3_420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val3_420_140_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val4_492_144_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val4_492_144_buf_req_0;
      n_fetch_val4_492_144_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val4_492_144_buf_req_1;
      n_fetch_val4_492_144_buf_ack_1<= rack(0);
      n_fetch_val4_492_144_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val4_492_144_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val4_492,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val4_492_144_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter_168_128_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter_168_128_buf_req_0;
      n_mycounter_168_128_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter_168_128_buf_req_1;
      n_mycounter_168_128_buf_ack_1<= rack(0);
      n_mycounter_168_128_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter_168_128_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter_168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter_168_128_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row1_186_149_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row1_186_149_buf_req_0;
      n_row1_186_149_buf_ack_0<= wack(0);
      rreq(0) <= n_row1_186_149_buf_req_1;
      n_row1_186_149_buf_ack_1<= rack(0);
      n_row1_186_149_buf : InterlockBuffer generic map ( -- 
        name => "n_row1_186_149_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row1_186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row1_186_149_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row2_194_154_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row2_194_154_buf_req_0;
      n_row2_194_154_buf_ack_0<= wack(0);
      rreq(0) <= n_row2_194_154_buf_req_1;
      n_row2_194_154_buf_ack_1<= rack(0);
      n_row2_194_154_buf : InterlockBuffer generic map ( -- 
        name => "n_row2_194_154_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row2_194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row2_194_154_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_110_inst_req_0;
      type_cast_110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_110_inst_req_1;
      type_cast_110_inst_ack_1<= rack(0);
      type_cast_110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_110_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_110_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_115_inst_req_0;
      type_cast_115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_115_inst_req_1;
      type_cast_115_inst_ack_1<= rack(0);
      type_cast_115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_115_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m2_factor_41,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_115_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_122_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_122_inst_req_0;
      type_cast_122_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_122_inst_req_1;
      type_cast_122_inst_ack_1<= rack(0);
      type_cast_122_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_122_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u32_u32_121_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_122_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_218_inst
    process(LSHR_u64_u64_217_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := LSHR_u64_u64_217_wire(7 downto 0);
      var_val1_219 <= tmp_var; -- 
    end process;
    type_cast_227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_227_inst_req_0;
      type_cast_227_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_227_inst_req_1;
      type_cast_227_inst_ack_1<= rack(0);
      type_cast_227_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_227_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_229_229_delayed_1_0_228,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_290_inst
    process(LSHR_u64_u64_289_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := LSHR_u64_u64_289_wire(7 downto 0);
      var_val2_291 <= tmp_var; -- 
    end process;
    type_cast_299_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_299_inst_req_0;
      type_cast_299_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_299_inst_req_1;
      type_cast_299_inst_ack_1<= rack(0);
      type_cast_299_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_299_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_289_289_delayed_1_0_300,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_35_inst
    process(MUL_u16_u16_34_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_34_wire(15 downto 0);
      m_factor_36 <= tmp_var; -- 
    end process;
    -- interlock type_cast_362_inst
    process(LSHR_u64_u64_361_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := LSHR_u64_u64_361_wire(7 downto 0);
      var_val3_363 <= tmp_var; -- 
    end process;
    type_cast_371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_371_inst_req_0;
      type_cast_371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_371_inst_req_1;
      type_cast_371_inst_ack_1<= rack(0);
      type_cast_371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_371_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_349_349_delayed_1_0_372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_434_inst
    process(LSHR_u64_u64_433_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := LSHR_u64_u64_433_wire(7 downto 0);
      var_val4_435 <= tmp_var; -- 
    end process;
    type_cast_443_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_443_inst_req_0;
      type_cast_443_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_443_inst_req_1;
      type_cast_443_inst_ack_1<= rack(0);
      type_cast_443_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_443_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_409_409_delayed_1_0_444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_60_inst
    process(LSHR_u32_u32_59_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_59_wire(31 downto 0);
      type_cast_60_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_74_inst
    process(LSHR_u32_u32_73_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_73_wire(31 downto 0);
      type_cast_74_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_92_inst
    process(ADD_u32_u32_91_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ADD_u32_u32_91_wire(31 downto 0);
      type_cast_92_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_254_index_1_rename
    process(LSHR_u64_u64_253_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_253_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_253_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_254_index_1_resize
    process(LSHR_u64_u64_253_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_253_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_253_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_254_root_address_inst
    process(array_obj_ref_254_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_254_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_254_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_326_index_1_rename
    process(LSHR_u64_u64_325_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_325_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_325_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_326_index_1_resize
    process(LSHR_u64_u64_325_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_325_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_325_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_326_root_address_inst
    process(array_obj_ref_326_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_326_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_326_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_index_1_rename
    process(LSHR_u64_u64_397_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_397_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_397_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_index_1_resize
    process(LSHR_u64_u64_397_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_397_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_397_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_root_address_inst
    process(array_obj_ref_398_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_398_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_398_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_470_index_1_rename
    process(LSHR_u64_u64_469_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_469_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_469_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_470_index_1_resize
    process(LSHR_u64_u64_469_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_469_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_469_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_470_root_address_inst
    process(array_obj_ref_470_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_470_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_470_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_index_1_rename
    process(type_cast_60_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_60_resized;
      ov(13 downto 0) := iv;
      type_cast_60_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_index_1_resize
    process(type_cast_60_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_60_wire;
      ov := iv(13 downto 0);
      type_cast_60_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_root_address_inst
    process(array_obj_ref_61_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_61_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_61_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_index_1_rename
    process(type_cast_74_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_74_resized;
      ov(13 downto 0) := iv;
      type_cast_74_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_index_1_resize
    process(type_cast_74_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_74_wire;
      ov := iv(13 downto 0);
      type_cast_74_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_root_address_inst
    process(array_obj_ref_75_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_75_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_75_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_93_index_1_rename
    process(type_cast_92_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_92_resized;
      ov(13 downto 0) := iv;
      type_cast_92_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_93_index_1_resize
    process(type_cast_92_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_92_wire;
      ov := iv(13 downto 0);
      type_cast_92_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_93_root_address_inst
    process(array_obj_ref_93_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_93_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_93_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_addr_0
    process(ptr_deref_263_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_263_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_263_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_base_resize
    process(fetch_addr1_256) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_256;
      ov := iv(13 downto 0);
      ptr_deref_263_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_gather_scatter
    process(ptr_deref_263_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_263_data_0;
      ov(63 downto 0) := iv;
      fv1_264 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_root_address_inst
    process(ptr_deref_263_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_263_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_263_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_335_addr_0
    process(ptr_deref_335_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_335_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_335_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_335_base_resize
    process(fetch_addr2_328) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_328;
      ov := iv(13 downto 0);
      ptr_deref_335_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_335_gather_scatter
    process(ptr_deref_335_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_335_data_0;
      ov(63 downto 0) := iv;
      fv2_336 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_335_root_address_inst
    process(ptr_deref_335_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_335_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_335_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_addr_0
    process(ptr_deref_407_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_407_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_407_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_base_resize
    process(fetch_addr3_400) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr3_400;
      ov := iv(13 downto 0);
      ptr_deref_407_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_gather_scatter
    process(ptr_deref_407_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_407_data_0;
      ov(63 downto 0) := iv;
      fv3_408 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_root_address_inst
    process(ptr_deref_407_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_407_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_407_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_addr_0
    process(ptr_deref_479_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_479_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_479_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_base_resize
    process(fetch_addr4_472) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr4_472;
      ov := iv(13 downto 0);
      ptr_deref_479_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_gather_scatter
    process(ptr_deref_479_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_479_data_0;
      ov(63 downto 0) := iv;
      fv4_480 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_root_address_inst
    process(ptr_deref_479_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_479_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_479_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_52_addr_0
    process(ptr_deref_52_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_52_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_52_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_52_base_resize
    process(fetch_add1_49) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add1_49;
      ov := iv(13 downto 0);
      ptr_deref_52_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_52_gather_scatter
    process(ptr_deref_52_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_52_data_0;
      ov(63 downto 0) := iv;
      my_fetch1_53 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_52_root_address_inst
    process(ptr_deref_52_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_52_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_52_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_addr_0
    process(ptr_deref_66_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_66_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_base_resize
    process(fetch_add2_63) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add2_63;
      ov := iv(13 downto 0);
      ptr_deref_66_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_gather_scatter
    process(ptr_deref_66_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_data_0;
      ov(63 downto 0) := iv;
      my_fetch2_67 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_root_address_inst
    process(ptr_deref_66_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_66_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_80_addr_0
    process(ptr_deref_80_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_80_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_80_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_80_base_resize
    process(fetch_add3_77) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add3_77;
      ov := iv(13 downto 0);
      ptr_deref_80_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_80_gather_scatter
    process(ptr_deref_80_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_80_data_0;
      ov(63 downto 0) := iv;
      my_fetch3_81 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_80_root_address_inst
    process(ptr_deref_80_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_80_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_80_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_98_addr_0
    process(ptr_deref_98_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_98_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_98_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_98_base_resize
    process(fetch_add4_95) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add4_95;
      ov := iv(13 downto 0);
      ptr_deref_98_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_98_gather_scatter
    process(ptr_deref_98_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_98_data_0;
      ov(63 downto 0) := iv;
      my_fetch4_99 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_98_root_address_inst
    process(ptr_deref_98_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_98_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_98_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_100_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue1_199;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_100_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_100_branch_req_0,
          ack0 => do_while_stmt_100_branch_ack_0,
          ack1 => do_while_stmt_100_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_183_inst
    process(row1_145) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row1_145, konst_182_wire_constant, tmp_var);
      ADD_u16_u16_183_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_191_inst
    process(row2_150) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row2_150, konst_190_wire_constant, tmp_var);
      ADD_u16_u16_191_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_121_inst
    process(m_factor_36, m2_factor_41) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, m2_factor_41, tmp_var);
      ADD_u32_u32_121_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_166_inst
    process(mycounter_124) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycounter_124, konst_165_wire_constant, tmp_var);
      ADD_u32_u32_166_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_91_inst
    process(LSHR_u32_u32_87_wire, LSHR_u32_u32_90_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(LSHR_u32_u32_87_wire, LSHR_u32_u32_90_wire, tmp_var);
      ADD_u32_u32_91_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_223_inst
    process(address1_102) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address1_102, konst_222_wire_constant, tmp_var);
      temp_address1_224 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_233_inst
    process(temp_address1_224, type_cast_229_229_delayed_1_0_228) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(temp_address1_224, type_cast_229_229_delayed_1_0_228, tmp_var);
      ADD_u64_u64_233_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_295_inst
    process(address2_107) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address2_107, konst_294_wire_constant, tmp_var);
      temp_address2_296 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_305_inst
    process(temp_address2_296, type_cast_289_289_delayed_1_0_300) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(temp_address2_296, type_cast_289_289_delayed_1_0_300, tmp_var);
      ADD_u64_u64_305_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_367_inst
    process(address3_112) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address3_112, konst_366_wire_constant, tmp_var);
      temp_address3_368 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_377_inst
    process(temp_address3_368, type_cast_349_349_delayed_1_0_372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(temp_address3_368, type_cast_349_349_delayed_1_0_372, tmp_var);
      ADD_u64_u64_377_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_439_inst
    process(address4_117) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address4_117, konst_438_wire_constant, tmp_var);
      temp_address4_440 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_449_inst
    process(temp_address4_440, type_cast_409_409_delayed_1_0_444) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(temp_address4_440, type_cast_409_409_delayed_1_0_444, tmp_var);
      ADD_u64_u64_449_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_246_inst
    process(NEQ_u64_u1_244_wire, continue1_199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_244_wire, continue1_199, tmp_var);
      fn1_247 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_318_inst
    process(NEQ_u64_u1_316_wire, continue1_199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_316_wire, continue1_199, tmp_var);
      fn2_319 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_390_inst
    process(NEQ_u64_u1_388_wire, continue1_199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_388_wire, continue1_199, tmp_var);
      fn3_391 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_462_inst
    process(NEQ_u64_u1_460_wire, continue2_204) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_460_wire, continue2_204, tmp_var);
      fn4_463 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_209_inst
    process(address1_102) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address1_102, konst_208_wire_constant, tmp_var);
      AND_u64_u64_209_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_281_inst
    process(address2_107) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address2_107, konst_280_wire_constant, tmp_var);
      AND_u64_u64_281_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_353_inst
    process(address3_112) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address3_112, konst_352_wire_constant, tmp_var);
      AND_u64_u64_353_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_425_inst
    process(address4_117) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address4_117, konst_424_wire_constant, tmp_var);
      AND_u64_u64_425_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_159_inst
    process(mycounter_124, m_factor_36) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycounter_124, m_factor_36, tmp_var);
      next_row_160 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_59_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_36, konst_58_wire_constant, tmp_var);
      LSHR_u32_u32_59_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_73_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_36, konst_72_wire_constant, tmp_var);
      LSHR_u32_u32_73_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_87_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_36, konst_86_wire_constant, tmp_var);
      LSHR_u32_u32_87_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_90_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_36, konst_89_wire_constant, tmp_var);
      LSHR_u32_u32_90_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_217_inst
    process(fetch_val1_129, my_num1_213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val1_129, my_num1_213, tmp_var);
      LSHR_u64_u64_217_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_240_inst
    process(n_address1_236) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address1_236, konst_239_wire_constant, tmp_var);
      LSHR_u64_u64_240_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_243_inst
    process(address1_102) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address1_102, konst_242_wire_constant, tmp_var);
      LSHR_u64_u64_243_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_253_inst
    process(n_address1_236) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address1_236, konst_252_wire_constant, tmp_var);
      LSHR_u64_u64_253_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_289_inst
    process(fetch_val2_133, my_num2_285) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val2_133, my_num2_285, tmp_var);
      LSHR_u64_u64_289_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_312_inst
    process(n_address2_308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address2_308, konst_311_wire_constant, tmp_var);
      LSHR_u64_u64_312_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_315_inst
    process(address2_107) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address2_107, konst_314_wire_constant, tmp_var);
      LSHR_u64_u64_315_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_325_inst
    process(n_address2_308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address2_308, konst_324_wire_constant, tmp_var);
      LSHR_u64_u64_325_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_361_inst
    process(fetch_val3_137, my_num3_357) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val3_137, my_num3_357, tmp_var);
      LSHR_u64_u64_361_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_384_inst
    process(n_address3_380) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address3_380, konst_383_wire_constant, tmp_var);
      LSHR_u64_u64_384_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_387_inst
    process(address3_112) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address3_112, konst_386_wire_constant, tmp_var);
      LSHR_u64_u64_387_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_397_inst
    process(n_address3_380) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address3_380, konst_396_wire_constant, tmp_var);
      LSHR_u64_u64_397_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_433_inst
    process(fetch_val4_141, my_num4_429) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val4_141, my_num4_429, tmp_var);
      LSHR_u64_u64_433_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_456_inst
    process(n_address4_452) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address4_452, konst_455_wire_constant, tmp_var);
      LSHR_u64_u64_456_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_459_inst
    process(address4_117) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address4_117, konst_458_wire_constant, tmp_var);
      LSHR_u64_u64_459_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_469_inst
    process(n_address4_452) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address4_452, konst_468_wire_constant, tmp_var);
      LSHR_u64_u64_469_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_34_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_34_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_244_inst
    process(LSHR_u64_u64_240_wire, LSHR_u64_u64_243_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_240_wire, LSHR_u64_u64_243_wire, tmp_var);
      NEQ_u64_u1_244_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_316_inst
    process(LSHR_u64_u64_312_wire, LSHR_u64_u64_315_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_312_wire, LSHR_u64_u64_315_wire, tmp_var);
      NEQ_u64_u1_316_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_388_inst
    process(LSHR_u64_u64_384_wire, LSHR_u64_u64_387_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_384_wire, LSHR_u64_u64_387_wire, tmp_var);
      NEQ_u64_u1_388_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_460_inst
    process(LSHR_u64_u64_456_wire, LSHR_u64_u64_459_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_456_wire, LSHR_u64_u64_459_wire, tmp_var);
      NEQ_u64_u1_460_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_40_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(m_factor_36, konst_39_wire_constant, tmp_var);
      m2_factor_41 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_212_inst
    process(SUB_u64_u64_210_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_210_wire, konst_211_wire_constant, tmp_var);
      my_num1_213 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_284_inst
    process(SUB_u64_u64_282_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_282_wire, konst_283_wire_constant, tmp_var);
      my_num2_285 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_356_inst
    process(SUB_u64_u64_354_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_354_wire, konst_355_wire_constant, tmp_var);
      my_num3_357 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_428_inst
    process(SUB_u64_u64_426_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_426_wire, konst_427_wire_constant, tmp_var);
      my_num4_429 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_210_inst
    process(konst_206_wire_constant, AND_u64_u64_209_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_206_wire_constant, AND_u64_u64_209_wire, tmp_var);
      SUB_u64_u64_210_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_282_inst
    process(konst_278_wire_constant, AND_u64_u64_281_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_278_wire_constant, AND_u64_u64_281_wire, tmp_var);
      SUB_u64_u64_282_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_354_inst
    process(konst_350_wire_constant, AND_u64_u64_353_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_350_wire_constant, AND_u64_u64_353_wire, tmp_var);
      SUB_u64_u64_354_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_426_inst
    process(konst_422_wire_constant, AND_u64_u64_425_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_422_wire_constant, AND_u64_u64_425_wire, tmp_var);
      SUB_u64_u64_426_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_172_inst
    process(row1_145, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row1_145, row_in_buffer, tmp_var);
      send_now1_173 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_177_inst
    process(row2_150, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row2_150, row_in_buffer, tmp_var);
      send_now2_178 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_198_inst
    process(n_row1_186, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row1_186, row_in_buffer, tmp_var);
      continue1_199 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_203_inst
    process(n_row2_194, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row2_194, row_in_buffer, tmp_var);
      continue2_204 <= tmp_var; --
    end process;
    -- shared split operator group (60) : array_obj_ref_254_index_offset 
    ApIntAdd_group_60: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_253_scaled;
      array_obj_ref_254_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_254_index_offset_req_0;
      array_obj_ref_254_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_254_index_offset_req_1;
      array_obj_ref_254_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_60_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_60_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_60",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : array_obj_ref_326_index_offset 
    ApIntAdd_group_61: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_325_scaled;
      array_obj_ref_326_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_326_index_offset_req_0;
      array_obj_ref_326_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_326_index_offset_req_1;
      array_obj_ref_326_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_61_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_61_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_61",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : array_obj_ref_398_index_offset 
    ApIntAdd_group_62: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_397_scaled;
      array_obj_ref_398_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_398_index_offset_req_0;
      array_obj_ref_398_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_398_index_offset_req_1;
      array_obj_ref_398_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_62_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_62_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_62",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : array_obj_ref_470_index_offset 
    ApIntAdd_group_63: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_469_scaled;
      array_obj_ref_470_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_470_index_offset_req_0;
      array_obj_ref_470_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_470_index_offset_req_1;
      array_obj_ref_470_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_63_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_63_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_63",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : array_obj_ref_61_index_offset 
    ApIntAdd_group_64: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_60_scaled;
      array_obj_ref_61_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_61_index_offset_req_0;
      array_obj_ref_61_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_61_index_offset_req_1;
      array_obj_ref_61_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_64_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_64_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_64",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : array_obj_ref_75_index_offset 
    ApIntAdd_group_65: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_74_scaled;
      array_obj_ref_75_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_75_index_offset_req_0;
      array_obj_ref_75_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_75_index_offset_req_1;
      array_obj_ref_75_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_65_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_65_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_65",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : array_obj_ref_93_index_offset 
    ApIntAdd_group_66: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_92_scaled;
      array_obj_ref_93_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_93_index_offset_req_0;
      array_obj_ref_93_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_93_index_offset_req_1;
      array_obj_ref_93_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_66_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_66_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_66",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared load operator group (0) : ptr_deref_52_load_0 ptr_deref_66_load_0 ptr_deref_407_load_0 ptr_deref_479_load_0 ptr_deref_80_load_0 ptr_deref_98_load_0 ptr_deref_263_load_0 ptr_deref_335_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(111 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 2, 4 => 2, 3 => 0, 2 => 0, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 2, 4 => 2, 3 => 1, 2 => 1, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => true, 1 => true, 2 => false, 3 => false, 4 => true, 5 => true, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 6, 1 => 6, 2 => 2, 3 => 2, 4 => 6, 5 => 6, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= ptr_deref_52_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_66_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_407_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_479_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_80_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_98_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_263_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_335_load_0_req_0;
      ptr_deref_52_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_66_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_407_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_479_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_80_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_98_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_263_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_335_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_52_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_66_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_407_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_479_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_80_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_98_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_263_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_335_load_0_req_1;
      ptr_deref_52_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_66_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_407_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_479_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_80_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_98_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_263_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_335_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn2_314_delayed_7_0_331(0);
      guard_vector(1)  <= fn1_254_delayed_7_0_259(0);
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <= fn4_434_delayed_7_0_475(0);
      guard_vector(5)  <= fn3_374_delayed_7_0_403(0);
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 2) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 2) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_52_word_address_0 & ptr_deref_66_word_address_0 & ptr_deref_407_word_address_0 & ptr_deref_479_word_address_0 & ptr_deref_80_word_address_0 & ptr_deref_98_word_address_0 & ptr_deref_263_word_address_0 & ptr_deref_335_word_address_0;
      ptr_deref_52_data_0 <= data_out(511 downto 448);
      ptr_deref_66_data_0 <= data_out(447 downto 384);
      ptr_deref_407_data_0 <= data_out(383 downto 320);
      ptr_deref_479_data_0 <= data_out(319 downto 256);
      ptr_deref_80_data_0 <= data_out(255 downto 192);
      ptr_deref_98_data_0 <= data_out(191 downto 128);
      ptr_deref_263_data_0 <= data_out(127 downto 64);
      ptr_deref_335_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_494_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe1_494_inst_req_0;
      WPIPE_input_pipe1_494_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe1_494_inst_req_1;
      WPIPE_input_pipe1_494_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_now1_173(0);
      data_in <= var_val1_219;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_input_pipe2_498_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe2_498_inst_req_0;
      WPIPE_input_pipe2_498_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe2_498_inst_req_1;
      WPIPE_input_pipe2_498_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_now1_173(0);
      data_in <= var_val2_291;
      input_pipe2_write_1_gI: SplitGuardInterface generic map(name => "input_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "input_pipe2", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe2_pipe_write_req(0),
          oack => input_pipe2_pipe_write_ack(0),
          odata => input_pipe2_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_input_pipe3_502_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe3_502_inst_req_0;
      WPIPE_input_pipe3_502_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe3_502_inst_req_1;
      WPIPE_input_pipe3_502_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_now1_173(0);
      data_in <= var_val3_363;
      input_pipe3_write_2_gI: SplitGuardInterface generic map(name => "input_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "input_pipe3", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe3_pipe_write_req(0),
          oack => input_pipe3_pipe_write_ack(0),
          odata => input_pipe3_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_input_pipe4_506_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe4_506_inst_req_0;
      WPIPE_input_pipe4_506_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe4_506_inst_req_1;
      WPIPE_input_pipe4_506_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_now2_178(0);
      data_in <= var_val4_435;
      input_pipe4_write_3_gI: SplitGuardInterface generic map(name => "input_pipe4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe4_write_3: OutputPortRevised -- 
        generic map ( name => "input_pipe4", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe4_pipe_write_req(0),
          oack => input_pipe4_pipe_write_ack(0),
          odata => input_pipe4_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(47 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(79 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    sendB_call_reqs : out  std_logic_vector(0 downto 0);
    sendB_call_acks : in   std_logic_vector(0 downto 0);
    sendB_call_data : out  std_logic_vector(31 downto 0);
    sendB_call_tag  :  out  std_logic_vector(0 downto 0);
    sendB_return_reqs : out  std_logic_vector(0 downto 0);
    sendB_return_acks : in   std_logic_vector(0 downto 0);
    sendB_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_3583_start: Boolean;
  signal convolution3D_CP_3583_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(7 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(7 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(7 downto 0);
      input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(7 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(7 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_1230_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1217_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1255_inst_req_0 : boolean;
  signal ptr_deref_1854_store_0_req_0 : boolean;
  signal type_cast_1246_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1255_inst_ack_0 : boolean;
  signal type_cast_1234_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1217_inst_req_0 : boolean;
  signal type_cast_1913_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1217_inst_req_1 : boolean;
  signal type_cast_1234_inst_req_1 : boolean;
  signal type_cast_1246_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1230_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1217_inst_ack_1 : boolean;
  signal type_cast_1284_inst_ack_1 : boolean;
  signal type_cast_1284_inst_req_1 : boolean;
  signal type_cast_1271_inst_ack_0 : boolean;
  signal type_cast_1221_inst_req_0 : boolean;
  signal type_cast_1284_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1242_inst_req_1 : boolean;
  signal type_cast_1221_inst_ack_0 : boolean;
  signal type_cast_1271_inst_req_0 : boolean;
  signal type_cast_1913_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1242_inst_ack_1 : boolean;
  signal type_cast_1246_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1255_inst_ack_1 : boolean;
  signal type_cast_1259_inst_ack_0 : boolean;
  signal type_cast_1821_inst_req_1 : boolean;
  signal type_cast_1869_inst_req_1 : boolean;
  signal type_cast_1271_inst_req_1 : boolean;
  signal type_cast_1234_inst_ack_0 : boolean;
  signal type_cast_1271_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_ack_1 : boolean;
  signal type_cast_1821_inst_ack_0 : boolean;
  signal type_cast_1821_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1230_inst_ack_0 : boolean;
  signal type_cast_1284_inst_req_0 : boolean;
  signal type_cast_1259_inst_req_1 : boolean;
  signal type_cast_1221_inst_req_1 : boolean;
  signal ptr_deref_1854_store_0_ack_0 : boolean;
  signal type_cast_1246_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1267_inst_ack_1 : boolean;
  signal type_cast_1869_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1267_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1267_inst_ack_0 : boolean;
  signal type_cast_1755_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1230_inst_req_1 : boolean;
  signal type_cast_1259_inst_ack_1 : boolean;
  signal type_cast_1234_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1267_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1255_inst_req_1 : boolean;
  signal type_cast_1221_inst_ack_1 : boolean;
  signal type_cast_1259_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1305_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1305_inst_ack_0 : boolean;
  signal type_cast_1745_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1242_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1292_inst_req_0 : boolean;
  signal type_cast_1821_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1292_inst_ack_0 : boolean;
  signal type_cast_1869_inst_req_0 : boolean;
  signal type_cast_1296_inst_req_1 : boolean;
  signal type_cast_1296_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1305_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1305_inst_ack_1 : boolean;
  signal type_cast_1745_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1292_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1292_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1280_inst_ack_0 : boolean;
  signal type_cast_1861_inst_ack_1 : boolean;
  signal type_cast_1861_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1317_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1317_inst_ack_0 : boolean;
  signal type_cast_1745_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1317_inst_req_1 : boolean;
  signal type_cast_1309_inst_req_0 : boolean;
  signal type_cast_1309_inst_ack_0 : boolean;
  signal type_cast_1309_inst_req_1 : boolean;
  signal type_cast_1309_inst_ack_1 : boolean;
  signal type_cast_1755_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1242_inst_req_0 : boolean;
  signal type_cast_1869_inst_ack_0 : boolean;
  signal type_cast_1296_inst_req_0 : boolean;
  signal type_cast_1334_inst_req_0 : boolean;
  signal addr_of_1851_final_reg_req_0 : boolean;
  signal type_cast_1334_inst_ack_0 : boolean;
  signal type_cast_1334_inst_req_1 : boolean;
  signal type_cast_1334_inst_ack_1 : boolean;
  signal type_cast_1783_inst_ack_1 : boolean;
  signal type_cast_1861_inst_ack_0 : boolean;
  signal type_cast_1861_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_ack_1 : boolean;
  signal type_cast_1783_inst_req_1 : boolean;
  signal type_cast_1321_inst_req_0 : boolean;
  signal addr_of_1851_final_reg_ack_1 : boolean;
  signal type_cast_1321_inst_ack_0 : boolean;
  signal type_cast_1321_inst_req_1 : boolean;
  signal addr_of_1851_final_reg_req_1 : boolean;
  signal type_cast_1321_inst_ack_1 : boolean;
  signal type_cast_1745_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1330_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1330_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1330_inst_req_1 : boolean;
  signal addr_of_1851_final_reg_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1330_inst_ack_1 : boolean;
  signal if_stmt_1807_branch_req_0 : boolean;
  signal type_cast_1296_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1317_inst_ack_1 : boolean;
  signal if_stmt_1807_branch_ack_0 : boolean;
  signal if_stmt_1807_branch_ack_1 : boolean;
  signal type_cast_1346_inst_req_0 : boolean;
  signal type_cast_1346_inst_ack_0 : boolean;
  signal type_cast_1346_inst_req_1 : boolean;
  signal type_cast_1346_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1355_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1355_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1355_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1355_inst_ack_1 : boolean;
  signal type_cast_1783_inst_ack_0 : boolean;
  signal type_cast_1783_inst_req_0 : boolean;
  signal type_cast_1359_inst_req_0 : boolean;
  signal type_cast_1359_inst_ack_0 : boolean;
  signal type_cast_1865_inst_ack_1 : boolean;
  signal type_cast_1359_inst_req_1 : boolean;
  signal type_cast_1359_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1367_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1367_inst_ack_0 : boolean;
  signal type_cast_1736_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1367_inst_req_1 : boolean;
  signal array_obj_ref_1850_index_offset_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1367_inst_ack_1 : boolean;
  signal if_stmt_1892_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1779_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1779_inst_req_1 : boolean;
  signal type_cast_1865_inst_req_1 : boolean;
  signal type_cast_1371_inst_req_0 : boolean;
  signal array_obj_ref_1850_index_offset_req_1 : boolean;
  signal type_cast_1371_inst_ack_0 : boolean;
  signal type_cast_1371_inst_req_1 : boolean;
  signal type_cast_1371_inst_ack_1 : boolean;
  signal type_cast_1736_inst_req_1 : boolean;
  signal type_cast_1913_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1380_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1380_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1380_inst_req_1 : boolean;
  signal array_obj_ref_1850_index_offset_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1380_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1779_inst_ack_0 : boolean;
  signal if_stmt_1892_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1779_inst_req_0 : boolean;
  signal type_cast_1384_inst_req_0 : boolean;
  signal array_obj_ref_1850_index_offset_req_0 : boolean;
  signal type_cast_1384_inst_ack_0 : boolean;
  signal type_cast_1865_inst_ack_0 : boolean;
  signal type_cast_1384_inst_req_1 : boolean;
  signal type_cast_1384_inst_ack_1 : boolean;
  signal type_cast_1736_inst_ack_0 : boolean;
  signal ptr_deref_1854_store_0_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_ack_0 : boolean;
  signal type_cast_1736_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1392_inst_ack_1 : boolean;
  signal type_cast_1759_inst_ack_1 : boolean;
  signal type_cast_1759_inst_req_1 : boolean;
  signal type_cast_1865_inst_req_0 : boolean;
  signal type_cast_1396_inst_req_0 : boolean;
  signal type_cast_1396_inst_ack_0 : boolean;
  signal type_cast_1396_inst_req_1 : boolean;
  signal type_cast_1396_inst_ack_1 : boolean;
  signal ptr_deref_1854_store_0_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_ack_1 : boolean;
  signal type_cast_1913_inst_req_0 : boolean;
  signal if_stmt_1892_branch_req_0 : boolean;
  signal type_cast_1759_inst_ack_0 : boolean;
  signal type_cast_1759_inst_req_0 : boolean;
  signal type_cast_1409_inst_req_0 : boolean;
  signal type_cast_1409_inst_ack_0 : boolean;
  signal type_cast_1409_inst_req_1 : boolean;
  signal type_cast_1409_inst_ack_1 : boolean;
  signal type_cast_1418_inst_req_0 : boolean;
  signal type_cast_1418_inst_ack_0 : boolean;
  signal type_cast_1418_inst_req_1 : boolean;
  signal type_cast_1418_inst_ack_1 : boolean;
  signal type_cast_1755_inst_ack_1 : boolean;
  signal type_cast_1755_inst_req_1 : boolean;
  signal if_stmt_1727_branch_ack_1 : boolean;
  signal type_cast_1422_inst_req_0 : boolean;
  signal type_cast_1422_inst_ack_0 : boolean;
  signal type_cast_1422_inst_req_1 : boolean;
  signal type_cast_1422_inst_ack_1 : boolean;
  signal if_stmt_1727_branch_ack_0 : boolean;
  signal WPIPE_output_pipe_2313_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2372_inst_ack_1 : boolean;
  signal if_stmt_1440_branch_req_0 : boolean;
  signal if_stmt_1440_branch_ack_1 : boolean;
  signal if_stmt_1440_branch_ack_0 : boolean;
  signal type_cast_1471_inst_req_0 : boolean;
  signal type_cast_1471_inst_ack_0 : boolean;
  signal type_cast_1471_inst_req_1 : boolean;
  signal type_cast_1471_inst_ack_1 : boolean;
  signal type_cast_2272_inst_req_1 : boolean;
  signal type_cast_2272_inst_ack_1 : boolean;
  signal type_cast_1480_inst_req_0 : boolean;
  signal type_cast_1480_inst_ack_0 : boolean;
  signal type_cast_1480_inst_req_1 : boolean;
  signal type_cast_1480_inst_ack_1 : boolean;
  signal addr_of_2302_final_reg_ack_1 : boolean;
  signal type_cast_1514_inst_req_0 : boolean;
  signal type_cast_1514_inst_ack_0 : boolean;
  signal type_cast_1514_inst_req_1 : boolean;
  signal type_cast_1514_inst_ack_1 : boolean;
  signal array_obj_ref_1536_index_offset_req_0 : boolean;
  signal array_obj_ref_1536_index_offset_ack_0 : boolean;
  signal array_obj_ref_1536_index_offset_req_1 : boolean;
  signal array_obj_ref_1536_index_offset_ack_1 : boolean;
  signal WPIPE_output_pipe_2316_inst_req_0 : boolean;
  signal WPIPE_output_pipe_2316_inst_ack_0 : boolean;
  signal type_cast_2441_inst_req_1 : boolean;
  signal addr_of_1537_final_reg_req_0 : boolean;
  signal addr_of_1537_final_reg_ack_0 : boolean;
  signal addr_of_1537_final_reg_req_1 : boolean;
  signal addr_of_1537_final_reg_ack_1 : boolean;
  signal if_stmt_2402_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1540_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1540_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1540_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1540_inst_ack_1 : boolean;
  signal array_obj_ref_2301_index_offset_req_0 : boolean;
  signal type_cast_2441_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2316_inst_req_1 : boolean;
  signal type_cast_1544_inst_req_0 : boolean;
  signal type_cast_1544_inst_ack_0 : boolean;
  signal type_cast_1544_inst_req_1 : boolean;
  signal type_cast_1544_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2316_inst_ack_1 : boolean;
  signal array_obj_ref_2301_index_offset_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1553_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1553_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1553_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1553_inst_ack_1 : boolean;
  signal call_stmt_2424_call_req_0 : boolean;
  signal type_cast_1557_inst_req_0 : boolean;
  signal type_cast_1557_inst_ack_0 : boolean;
  signal type_cast_1557_inst_req_1 : boolean;
  signal type_cast_1557_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1571_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1571_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1571_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1571_inst_ack_1 : boolean;
  signal if_stmt_2402_branch_ack_1 : boolean;
  signal WPIPE_output_pipe_2319_inst_req_0 : boolean;
  signal type_cast_1575_inst_req_0 : boolean;
  signal type_cast_1575_inst_ack_0 : boolean;
  signal type_cast_1575_inst_req_1 : boolean;
  signal type_cast_1575_inst_ack_1 : boolean;
  signal type_cast_2458_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_2375_inst_req_0 : boolean;
  signal WPIPE_output_pipe_2319_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1589_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1589_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1589_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1589_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2319_inst_req_1 : boolean;
  signal WPIPE_output_pipe_2319_inst_ack_1 : boolean;
  signal call_stmt_2424_call_ack_0 : boolean;
  signal type_cast_1593_inst_req_0 : boolean;
  signal type_cast_1593_inst_ack_0 : boolean;
  signal type_cast_1593_inst_req_1 : boolean;
  signal type_cast_1593_inst_ack_1 : boolean;
  signal array_obj_ref_2301_index_offset_req_1 : boolean;
  signal type_cast_2413_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1607_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1607_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1607_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1607_inst_ack_1 : boolean;
  signal type_cast_2413_inst_ack_0 : boolean;
  signal type_cast_1611_inst_req_0 : boolean;
  signal type_cast_1611_inst_ack_0 : boolean;
  signal type_cast_1611_inst_req_1 : boolean;
  signal type_cast_1611_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1625_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1625_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1625_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1625_inst_ack_1 : boolean;
  signal type_cast_1629_inst_req_0 : boolean;
  signal type_cast_1629_inst_ack_0 : boolean;
  signal type_cast_1629_inst_req_1 : boolean;
  signal type_cast_1629_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1643_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1643_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1643_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1643_inst_ack_1 : boolean;
  signal type_cast_1647_inst_req_0 : boolean;
  signal type_cast_1647_inst_ack_0 : boolean;
  signal type_cast_1647_inst_req_1 : boolean;
  signal type_cast_1647_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1661_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1661_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1661_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1661_inst_ack_1 : boolean;
  signal type_cast_1665_inst_req_0 : boolean;
  signal type_cast_1665_inst_ack_0 : boolean;
  signal type_cast_1665_inst_req_1 : boolean;
  signal type_cast_1665_inst_ack_1 : boolean;
  signal ptr_deref_1673_store_0_req_0 : boolean;
  signal ptr_deref_1673_store_0_ack_0 : boolean;
  signal ptr_deref_1673_store_0_req_1 : boolean;
  signal ptr_deref_1673_store_0_ack_1 : boolean;
  signal if_stmt_1687_branch_req_0 : boolean;
  signal if_stmt_1687_branch_ack_1 : boolean;
  signal if_stmt_1687_branch_ack_0 : boolean;
  signal type_cast_1703_inst_req_0 : boolean;
  signal type_cast_1703_inst_ack_0 : boolean;
  signal type_cast_1703_inst_req_1 : boolean;
  signal type_cast_1703_inst_ack_1 : boolean;
  signal if_stmt_1727_branch_req_0 : boolean;
  signal type_cast_1917_inst_req_0 : boolean;
  signal type_cast_1917_inst_ack_0 : boolean;
  signal type_cast_1917_inst_req_1 : boolean;
  signal type_cast_1917_inst_ack_1 : boolean;
  signal type_cast_1926_inst_req_0 : boolean;
  signal type_cast_1926_inst_ack_0 : boolean;
  signal type_cast_1926_inst_req_1 : boolean;
  signal type_cast_1926_inst_ack_1 : boolean;
  signal type_cast_1935_inst_req_0 : boolean;
  signal type_cast_1935_inst_ack_0 : boolean;
  signal type_cast_1935_inst_req_1 : boolean;
  signal type_cast_1935_inst_ack_1 : boolean;
  signal type_cast_1969_inst_req_0 : boolean;
  signal type_cast_1969_inst_ack_0 : boolean;
  signal type_cast_1969_inst_req_1 : boolean;
  signal type_cast_1969_inst_ack_1 : boolean;
  signal addr_of_2302_final_reg_req_1 : boolean;
  signal WPIPE_output_pipe_2313_inst_req_1 : boolean;
  signal array_obj_ref_1991_index_offset_req_0 : boolean;
  signal WPIPE_num_out_pipe_2372_inst_req_1 : boolean;
  signal array_obj_ref_1991_index_offset_ack_0 : boolean;
  signal array_obj_ref_1991_index_offset_req_1 : boolean;
  signal array_obj_ref_1991_index_offset_ack_1 : boolean;
  signal type_cast_2441_inst_ack_0 : boolean;
  signal type_cast_2441_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_2372_inst_ack_0 : boolean;
  signal addr_of_1992_final_reg_req_0 : boolean;
  signal WPIPE_num_out_pipe_2372_inst_req_0 : boolean;
  signal addr_of_1992_final_reg_ack_0 : boolean;
  signal addr_of_1992_final_reg_req_1 : boolean;
  signal addr_of_1992_final_reg_ack_1 : boolean;
  signal WPIPE_output_pipe_2313_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_2313_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1995_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1995_inst_ack_0 : boolean;
  signal addr_of_2302_final_reg_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1995_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1995_inst_ack_1 : boolean;
  signal call_stmt_2390_call_ack_1 : boolean;
  signal RPIPE_input_done_pipe_2420_inst_ack_1 : boolean;
  signal type_cast_1999_inst_req_0 : boolean;
  signal type_cast_1999_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2420_inst_req_1 : boolean;
  signal type_cast_1999_inst_req_1 : boolean;
  signal type_cast_1999_inst_ack_1 : boolean;
  signal call_stmt_2390_call_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2008_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2008_inst_ack_0 : boolean;
  signal addr_of_2302_final_reg_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2008_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2008_inst_ack_1 : boolean;
  signal type_cast_2437_inst_ack_1 : boolean;
  signal type_cast_2437_inst_req_1 : boolean;
  signal type_cast_2012_inst_req_0 : boolean;
  signal type_cast_2012_inst_ack_0 : boolean;
  signal type_cast_2012_inst_req_1 : boolean;
  signal type_cast_2350_inst_ack_1 : boolean;
  signal type_cast_2012_inst_ack_1 : boolean;
  signal type_cast_2468_inst_ack_0 : boolean;
  signal type_cast_2468_inst_ack_1 : boolean;
  signal call_stmt_2390_call_ack_0 : boolean;
  signal call_stmt_2312_call_ack_1 : boolean;
  signal call_stmt_2312_call_req_1 : boolean;
  signal type_cast_2350_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2026_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2026_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2026_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2026_inst_ack_1 : boolean;
  signal type_cast_2030_inst_req_0 : boolean;
  signal type_cast_2030_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2420_inst_ack_0 : boolean;
  signal type_cast_2030_inst_req_1 : boolean;
  signal type_cast_2350_inst_ack_0 : boolean;
  signal type_cast_2030_inst_ack_1 : boolean;
  signal type_cast_2468_inst_req_0 : boolean;
  signal call_stmt_2454_call_ack_1 : boolean;
  signal type_cast_2468_inst_req_1 : boolean;
  signal call_stmt_2454_call_req_1 : boolean;
  signal call_stmt_2390_call_req_0 : boolean;
  signal call_stmt_2312_call_ack_0 : boolean;
  signal call_stmt_2312_call_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2044_inst_req_0 : boolean;
  signal type_cast_2350_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2044_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2044_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2044_inst_ack_1 : boolean;
  signal type_cast_2437_inst_ack_0 : boolean;
  signal type_cast_2437_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_2420_inst_req_0 : boolean;
  signal type_cast_2048_inst_req_0 : boolean;
  signal type_cast_2048_inst_ack_0 : boolean;
  signal type_cast_2048_inst_req_1 : boolean;
  signal type_cast_2048_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2062_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2062_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2062_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2062_inst_ack_1 : boolean;
  signal type_cast_2458_inst_ack_1 : boolean;
  signal type_cast_2428_inst_ack_1 : boolean;
  signal type_cast_2428_inst_req_1 : boolean;
  signal type_cast_2066_inst_req_0 : boolean;
  signal type_cast_2341_inst_ack_1 : boolean;
  signal type_cast_2066_inst_ack_0 : boolean;
  signal type_cast_2066_inst_req_1 : boolean;
  signal type_cast_2341_inst_req_1 : boolean;
  signal type_cast_2066_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2080_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2080_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2080_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2080_inst_ack_1 : boolean;
  signal type_cast_2458_inst_req_1 : boolean;
  signal type_cast_2428_inst_ack_0 : boolean;
  signal type_cast_2428_inst_req_0 : boolean;
  signal call_stmt_2386_call_ack_1 : boolean;
  signal ptr_deref_2305_store_0_ack_1 : boolean;
  signal type_cast_2084_inst_req_0 : boolean;
  signal type_cast_2341_inst_ack_0 : boolean;
  signal type_cast_2084_inst_ack_0 : boolean;
  signal type_cast_2084_inst_req_1 : boolean;
  signal type_cast_2341_inst_req_0 : boolean;
  signal type_cast_2084_inst_ack_1 : boolean;
  signal call_stmt_2454_call_ack_0 : boolean;
  signal call_stmt_2454_call_req_0 : boolean;
  signal call_stmt_2386_call_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2098_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2098_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2098_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2098_inst_ack_1 : boolean;
  signal ptr_deref_2305_store_0_req_1 : boolean;
  signal call_stmt_2386_call_ack_0 : boolean;
  signal type_cast_2102_inst_req_0 : boolean;
  signal type_cast_2102_inst_ack_0 : boolean;
  signal type_cast_2102_inst_req_1 : boolean;
  signal type_cast_2102_inst_ack_1 : boolean;
  signal call_stmt_2386_call_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2116_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2116_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2116_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2116_inst_ack_1 : boolean;
  signal type_cast_2413_inst_ack_1 : boolean;
  signal type_cast_2120_inst_req_0 : boolean;
  signal type_cast_2331_inst_ack_1 : boolean;
  signal type_cast_2120_inst_ack_0 : boolean;
  signal type_cast_2120_inst_req_1 : boolean;
  signal type_cast_2331_inst_req_1 : boolean;
  signal type_cast_2120_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2375_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2375_inst_req_1 : boolean;
  signal type_cast_2331_inst_ack_0 : boolean;
  signal if_stmt_2402_branch_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2416_inst_ack_1 : boolean;
  signal type_cast_2331_inst_req_0 : boolean;
  signal ptr_deref_2128_store_0_req_0 : boolean;
  signal ptr_deref_2305_store_0_ack_0 : boolean;
  signal ptr_deref_2128_store_0_ack_0 : boolean;
  signal type_cast_2272_inst_ack_0 : boolean;
  signal ptr_deref_2128_store_0_req_1 : boolean;
  signal ptr_deref_2305_store_0_req_0 : boolean;
  signal ptr_deref_2128_store_0_ack_1 : boolean;
  signal type_cast_2458_inst_ack_0 : boolean;
  signal type_cast_2413_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_2416_inst_req_1 : boolean;
  signal type_cast_2272_inst_req_0 : boolean;
  signal if_stmt_2142_branch_req_0 : boolean;
  signal if_stmt_2142_branch_ack_1 : boolean;
  signal if_stmt_2142_branch_ack_0 : boolean;
  signal type_cast_2158_inst_req_0 : boolean;
  signal type_cast_2158_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2416_inst_ack_0 : boolean;
  signal type_cast_2158_inst_req_1 : boolean;
  signal type_cast_2158_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2375_inst_ack_0 : boolean;
  signal call_stmt_2424_call_ack_1 : boolean;
  signal call_stmt_2424_call_req_1 : boolean;
  signal RPIPE_input_done_pipe_2416_inst_req_0 : boolean;
  signal array_obj_ref_2301_index_offset_ack_1 : boolean;
  signal if_stmt_2182_branch_req_0 : boolean;
  signal if_stmt_2182_branch_ack_1 : boolean;
  signal if_stmt_2182_branch_ack_0 : boolean;
  signal type_cast_2206_inst_req_0 : boolean;
  signal type_cast_2206_inst_ack_0 : boolean;
  signal type_cast_2206_inst_req_1 : boolean;
  signal type_cast_2206_inst_ack_1 : boolean;
  signal type_cast_2210_inst_req_0 : boolean;
  signal type_cast_2210_inst_ack_0 : boolean;
  signal type_cast_2210_inst_req_1 : boolean;
  signal type_cast_2210_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2230_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2230_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2230_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2230_inst_ack_1 : boolean;
  signal type_cast_2234_inst_req_0 : boolean;
  signal type_cast_2234_inst_ack_0 : boolean;
  signal type_cast_2234_inst_req_1 : boolean;
  signal type_cast_2234_inst_ack_1 : boolean;
  signal if_stmt_2258_branch_req_0 : boolean;
  signal if_stmt_2258_branch_ack_1 : boolean;
  signal if_stmt_2258_branch_ack_0 : boolean;
  signal type_cast_2478_inst_req_0 : boolean;
  signal type_cast_2478_inst_ack_0 : boolean;
  signal type_cast_2478_inst_req_1 : boolean;
  signal type_cast_2478_inst_ack_1 : boolean;
  signal type_cast_2488_inst_req_0 : boolean;
  signal type_cast_2488_inst_ack_0 : boolean;
  signal type_cast_2488_inst_req_1 : boolean;
  signal type_cast_2488_inst_ack_1 : boolean;
  signal type_cast_2498_inst_req_0 : boolean;
  signal type_cast_2498_inst_ack_0 : boolean;
  signal type_cast_2498_inst_req_1 : boolean;
  signal type_cast_2498_inst_ack_1 : boolean;
  signal type_cast_2508_inst_req_0 : boolean;
  signal type_cast_2508_inst_ack_0 : boolean;
  signal type_cast_2508_inst_req_1 : boolean;
  signal type_cast_2508_inst_ack_1 : boolean;
  signal type_cast_2518_inst_req_0 : boolean;
  signal type_cast_2518_inst_ack_0 : boolean;
  signal type_cast_2518_inst_req_1 : boolean;
  signal type_cast_2518_inst_ack_1 : boolean;
  signal type_cast_2528_inst_req_0 : boolean;
  signal type_cast_2528_inst_ack_0 : boolean;
  signal type_cast_2528_inst_req_1 : boolean;
  signal type_cast_2528_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2530_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2530_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2530_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2530_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2533_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2533_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2533_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2533_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2536_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2536_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2536_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2536_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2539_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2539_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2539_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2539_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2542_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2542_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2542_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2542_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2545_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2545_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2545_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2545_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2548_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2548_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2548_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2548_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2551_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2551_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2551_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2551_inst_ack_1 : boolean;
  signal phi_stmt_1524_req_0 : boolean;
  signal type_cast_1530_inst_req_0 : boolean;
  signal type_cast_1530_inst_ack_0 : boolean;
  signal type_cast_1530_inst_req_1 : boolean;
  signal type_cast_1530_inst_ack_1 : boolean;
  signal phi_stmt_1524_req_1 : boolean;
  signal phi_stmt_1524_ack_0 : boolean;
  signal phi_stmt_1707_req_1 : boolean;
  signal type_cast_1710_inst_req_0 : boolean;
  signal type_cast_1710_inst_ack_0 : boolean;
  signal type_cast_1710_inst_req_1 : boolean;
  signal type_cast_1710_inst_ack_1 : boolean;
  signal phi_stmt_1707_req_0 : boolean;
  signal phi_stmt_1707_ack_0 : boolean;
  signal type_cast_1773_inst_req_0 : boolean;
  signal type_cast_1773_inst_ack_0 : boolean;
  signal type_cast_1773_inst_req_1 : boolean;
  signal type_cast_1773_inst_ack_1 : boolean;
  signal phi_stmt_1770_req_0 : boolean;
  signal type_cast_1766_inst_req_0 : boolean;
  signal type_cast_1766_inst_ack_0 : boolean;
  signal type_cast_1766_inst_req_1 : boolean;
  signal type_cast_1766_inst_ack_1 : boolean;
  signal phi_stmt_1763_req_0 : boolean;
  signal phi_stmt_1770_req_1 : boolean;
  signal phi_stmt_1763_req_1 : boolean;
  signal phi_stmt_1763_ack_0 : boolean;
  signal phi_stmt_1770_ack_0 : boolean;
  signal type_cast_1817_inst_req_0 : boolean;
  signal type_cast_1817_inst_ack_0 : boolean;
  signal type_cast_1817_inst_req_1 : boolean;
  signal type_cast_1817_inst_ack_1 : boolean;
  signal phi_stmt_1814_req_0 : boolean;
  signal phi_stmt_2359_ack_0 : boolean;
  signal phi_stmt_1814_ack_0 : boolean;
  signal phi_stmt_1979_req_0 : boolean;
  signal type_cast_1985_inst_req_0 : boolean;
  signal type_cast_1985_inst_ack_0 : boolean;
  signal type_cast_1985_inst_req_1 : boolean;
  signal type_cast_1985_inst_ack_1 : boolean;
  signal phi_stmt_1979_req_1 : boolean;
  signal phi_stmt_1979_ack_0 : boolean;
  signal type_cast_2165_inst_req_0 : boolean;
  signal type_cast_2165_inst_ack_0 : boolean;
  signal type_cast_2165_inst_req_1 : boolean;
  signal type_cast_2165_inst_ack_1 : boolean;
  signal phi_stmt_2162_req_0 : boolean;
  signal phi_stmt_2162_req_1 : boolean;
  signal phi_stmt_2162_ack_0 : boolean;
  signal type_cast_2227_inst_req_0 : boolean;
  signal type_cast_2227_inst_ack_0 : boolean;
  signal type_cast_2227_inst_req_1 : boolean;
  signal type_cast_2227_inst_ack_1 : boolean;
  signal phi_stmt_2221_req_1 : boolean;
  signal type_cast_2220_inst_req_0 : boolean;
  signal type_cast_2220_inst_ack_0 : boolean;
  signal type_cast_2220_inst_req_1 : boolean;
  signal type_cast_2220_inst_ack_1 : boolean;
  signal phi_stmt_2214_req_1 : boolean;
  signal phi_stmt_2221_req_0 : boolean;
  signal phi_stmt_2214_req_0 : boolean;
  signal phi_stmt_2214_ack_0 : boolean;
  signal phi_stmt_2221_ack_0 : boolean;
  signal type_cast_2268_inst_req_0 : boolean;
  signal type_cast_2268_inst_ack_0 : boolean;
  signal type_cast_2268_inst_req_1 : boolean;
  signal type_cast_2268_inst_ack_1 : boolean;
  signal phi_stmt_2265_req_0 : boolean;
  signal phi_stmt_2265_ack_0 : boolean;
  signal phi_stmt_2359_req_0 : boolean;
  signal type_cast_2365_inst_req_0 : boolean;
  signal type_cast_2365_inst_ack_0 : boolean;
  signal type_cast_2365_inst_req_1 : boolean;
  signal type_cast_2365_inst_ack_1 : boolean;
  signal phi_stmt_2359_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_3583_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_3583_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_3583_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_3583_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_3583: Block -- control-path 
    signal convolution3D_CP_3583_elements: BooleanArray(390 downto 0);
    -- 
  begin -- 
    convolution3D_CP_3583_elements(0) <= convolution3D_CP_3583_start;
    convolution3D_CP_3583_symbol <= convolution3D_CP_3583_elements(322);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0:  members (62) 
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1215/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439__entry__
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/branch_block_stmt_1215__entry__
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_Update/cr
      -- 
    rr_3703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => RPIPE_maxpool_input_pipe_1217_inst_req_0); -- 
    cr_3750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1234_inst_req_1); -- 
    cr_3778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1246_inst_req_1); -- 
    cr_3862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1284_inst_req_1); -- 
    cr_3834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1271_inst_req_1); -- 
    cr_3806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1259_inst_req_1); -- 
    cr_3722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1221_inst_req_1); -- 
    cr_3890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1296_inst_req_1); -- 
    cr_3918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1309_inst_req_1); -- 
    cr_3974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1334_inst_req_1); -- 
    cr_3946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1321_inst_req_1); -- 
    cr_4002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1346_inst_req_1); -- 
    cr_4030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1359_inst_req_1); -- 
    cr_4058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1371_inst_req_1); -- 
    cr_4086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1384_inst_req_1); -- 
    cr_4114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1396_inst_req_1); -- 
    cr_4142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1409_inst_req_1); -- 
    cr_4156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1418_inst_req_1); -- 
    cr_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(0), ack => type_cast_1422_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_update_start_
      -- 
    ra_3704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1217_inst_ack_0, ack => convolution3D_CP_3583_elements(1)); -- 
    cr_3708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(1), ack => RPIPE_maxpool_input_pipe_1217_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1217_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_sample_start_
      -- 
    ca_3709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1217_inst_ack_1, ack => convolution3D_CP_3583_elements(2)); -- 
    rr_3717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(2), ack => type_cast_1221_inst_req_0); -- 
    rr_3731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(2), ack => RPIPE_maxpool_input_pipe_1230_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_sample_completed_
      -- 
    ra_3718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_0, ack => convolution3D_CP_3583_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1221_update_completed_
      -- 
    ca_3723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_1, ack => convolution3D_CP_3583_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_Update/cr
      -- 
    ra_3732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1230_inst_ack_0, ack => convolution3D_CP_3583_elements(5)); -- 
    cr_3736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(5), ack => RPIPE_maxpool_input_pipe_1230_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1230_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_Sample/$entry
      -- 
    ca_3737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1230_inst_ack_1, ack => convolution3D_CP_3583_elements(6)); -- 
    rr_3745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(6), ack => type_cast_1234_inst_req_0); -- 
    rr_3759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(6), ack => RPIPE_maxpool_input_pipe_1242_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_Sample/$exit
      -- 
    ra_3746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_0, ack => convolution3D_CP_3583_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1234_Update/ca
      -- 
    ca_3751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_1, ack => convolution3D_CP_3583_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_Sample/$exit
      -- 
    ra_3760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1242_inst_ack_0, ack => convolution3D_CP_3583_elements(9)); -- 
    cr_3764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(9), ack => RPIPE_maxpool_input_pipe_1242_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1242_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_Sample/$entry
      -- 
    ca_3765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1242_inst_ack_1, ack => convolution3D_CP_3583_elements(10)); -- 
    rr_3773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(10), ack => type_cast_1246_inst_req_0); -- 
    rr_3787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(10), ack => RPIPE_maxpool_input_pipe_1255_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_Sample/$exit
      -- 
    ra_3774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1246_inst_ack_0, ack => convolution3D_CP_3583_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1246_Update/$exit
      -- 
    ca_3779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1246_inst_ack_1, ack => convolution3D_CP_3583_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_Update/cr
      -- 
    ra_3788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1255_inst_ack_0, ack => convolution3D_CP_3583_elements(13)); -- 
    cr_3792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(13), ack => RPIPE_maxpool_input_pipe_1255_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1255_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_sample_start_
      -- 
    ca_3793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1255_inst_ack_1, ack => convolution3D_CP_3583_elements(14)); -- 
    rr_3815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(14), ack => RPIPE_maxpool_input_pipe_1267_inst_req_0); -- 
    rr_3801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(14), ack => type_cast_1259_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_Sample/$exit
      -- 
    ra_3802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1259_inst_ack_0, ack => convolution3D_CP_3583_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1259_update_completed_
      -- 
    ca_3807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1259_inst_ack_1, ack => convolution3D_CP_3583_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_Update/cr
      -- 
    ra_3816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1267_inst_ack_0, ack => convolution3D_CP_3583_elements(17)); -- 
    cr_3820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(17), ack => RPIPE_maxpool_input_pipe_1267_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1267_Update/$exit
      -- 
    ca_3821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1267_inst_ack_1, ack => convolution3D_CP_3583_elements(18)); -- 
    rr_3843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(18), ack => RPIPE_maxpool_input_pipe_1280_inst_req_0); -- 
    rr_3829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(18), ack => type_cast_1271_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_sample_completed_
      -- 
    ra_3830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1271_inst_ack_0, ack => convolution3D_CP_3583_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1271_update_completed_
      -- 
    ca_3835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1271_inst_ack_1, ack => convolution3D_CP_3583_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_update_start_
      -- 
    ra_3844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1280_inst_ack_0, ack => convolution3D_CP_3583_elements(21)); -- 
    cr_3848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(21), ack => RPIPE_maxpool_input_pipe_1280_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1280_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_Sample/rr
      -- 
    ca_3849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1280_inst_ack_1, ack => convolution3D_CP_3583_elements(22)); -- 
    rr_3857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(22), ack => type_cast_1284_inst_req_0); -- 
    rr_3871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(22), ack => RPIPE_maxpool_input_pipe_1292_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_Sample/$exit
      -- 
    ra_3858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_0, ack => convolution3D_CP_3583_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1284_update_completed_
      -- 
    ca_3863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_1, ack => convolution3D_CP_3583_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_Update/$entry
      -- 
    ra_3872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1292_inst_ack_0, ack => convolution3D_CP_3583_elements(25)); -- 
    cr_3876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(25), ack => RPIPE_maxpool_input_pipe_1292_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1292_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_sample_start_
      -- 
    ca_3877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1292_inst_ack_1, ack => convolution3D_CP_3583_elements(26)); -- 
    rr_3885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(26), ack => type_cast_1296_inst_req_0); -- 
    rr_3899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(26), ack => RPIPE_maxpool_input_pipe_1305_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_Sample/ra
      -- 
    ra_3886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1296_inst_ack_0, ack => convolution3D_CP_3583_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	71 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1296_update_completed_
      -- 
    ca_3891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1296_inst_ack_1, ack => convolution3D_CP_3583_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_Update/cr
      -- CP-element group 29: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_update_start_
      -- 
    ra_3900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1305_inst_ack_0, ack => convolution3D_CP_3583_elements(29)); -- 
    cr_3904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(29), ack => RPIPE_maxpool_input_pipe_1305_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1305_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_Sample/$entry
      -- 
    ca_3905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1305_inst_ack_1, ack => convolution3D_CP_3583_elements(30)); -- 
    rr_3913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(30), ack => type_cast_1309_inst_req_0); -- 
    rr_3927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(30), ack => RPIPE_maxpool_input_pipe_1317_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_Sample/$exit
      -- 
    ra_3914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1309_inst_ack_0, ack => convolution3D_CP_3583_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	71 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1309_update_completed_
      -- 
    ca_3919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1309_inst_ack_1, ack => convolution3D_CP_3583_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_update_start_
      -- CP-element group 33: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_Update/cr
      -- 
    ra_3928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1317_inst_ack_0, ack => convolution3D_CP_3583_elements(33)); -- 
    cr_3932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(33), ack => RPIPE_maxpool_input_pipe_1317_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1317_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_sample_start_
      -- 
    ca_3933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1317_inst_ack_1, ack => convolution3D_CP_3583_elements(34)); -- 
    rr_3941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(34), ack => type_cast_1321_inst_req_0); -- 
    rr_3955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(34), ack => RPIPE_maxpool_input_pipe_1330_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_sample_completed_
      -- 
    ra_3942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1321_inst_ack_0, ack => convolution3D_CP_3583_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	71 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1321_update_completed_
      -- 
    ca_3947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1321_inst_ack_1, ack => convolution3D_CP_3583_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_Update/cr
      -- 
    ra_3956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1330_inst_ack_0, ack => convolution3D_CP_3583_elements(37)); -- 
    cr_3960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(37), ack => RPIPE_maxpool_input_pipe_1330_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1330_Update/ca
      -- 
    ca_3961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1330_inst_ack_1, ack => convolution3D_CP_3583_elements(38)); -- 
    rr_3969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(38), ack => type_cast_1334_inst_req_0); -- 
    rr_3983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(38), ack => RPIPE_maxpool_input_pipe_1342_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_Sample/ra
      -- 
    ra_3970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1334_inst_ack_0, ack => convolution3D_CP_3583_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	71 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1334_Update/ca
      -- 
    ca_3975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1334_inst_ack_1, ack => convolution3D_CP_3583_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_Update/cr
      -- 
    ra_3984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1342_inst_ack_0, ack => convolution3D_CP_3583_elements(41)); -- 
    cr_3988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(41), ack => RPIPE_maxpool_input_pipe_1342_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1342_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_Sample/rr
      -- 
    ca_3989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1342_inst_ack_1, ack => convolution3D_CP_3583_elements(42)); -- 
    rr_3997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(42), ack => type_cast_1346_inst_req_0); -- 
    rr_4011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(42), ack => RPIPE_maxpool_input_pipe_1355_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_Sample/ra
      -- 
    ra_3998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_0, ack => convolution3D_CP_3583_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	71 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1346_Update/ca
      -- 
    ca_4003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_1, ack => convolution3D_CP_3583_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_update_start_
      -- CP-element group 45: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_Update/cr
      -- 
    ra_4012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1355_inst_ack_0, ack => convolution3D_CP_3583_elements(45)); -- 
    cr_4016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(45), ack => RPIPE_maxpool_input_pipe_1355_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1355_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_Sample/rr
      -- 
    ca_4017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1355_inst_ack_1, ack => convolution3D_CP_3583_elements(46)); -- 
    rr_4025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(46), ack => type_cast_1359_inst_req_0); -- 
    rr_4039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(46), ack => RPIPE_maxpool_input_pipe_1367_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_Sample/ra
      -- 
    ra_4026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1359_inst_ack_0, ack => convolution3D_CP_3583_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	71 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1359_Update/ca
      -- 
    ca_4031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1359_inst_ack_1, ack => convolution3D_CP_3583_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_Update/cr
      -- 
    ra_4040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1367_inst_ack_0, ack => convolution3D_CP_3583_elements(49)); -- 
    cr_4044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(49), ack => RPIPE_maxpool_input_pipe_1367_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1367_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_Sample/rr
      -- 
    ca_4045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1367_inst_ack_1, ack => convolution3D_CP_3583_elements(50)); -- 
    rr_4053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(50), ack => type_cast_1371_inst_req_0); -- 
    rr_4067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(50), ack => RPIPE_maxpool_input_pipe_1380_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_Sample/ra
      -- 
    ra_4054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1371_inst_ack_0, ack => convolution3D_CP_3583_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	71 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1371_Update/ca
      -- 
    ca_4059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1371_inst_ack_1, ack => convolution3D_CP_3583_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_Update/cr
      -- 
    ra_4068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1380_inst_ack_0, ack => convolution3D_CP_3583_elements(53)); -- 
    cr_4072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(53), ack => RPIPE_maxpool_input_pipe_1380_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1380_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_Sample/rr
      -- 
    ca_4073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1380_inst_ack_1, ack => convolution3D_CP_3583_elements(54)); -- 
    rr_4095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(54), ack => RPIPE_maxpool_input_pipe_1392_inst_req_0); -- 
    rr_4081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(54), ack => type_cast_1384_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_Sample/ra
      -- 
    ra_4082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1384_inst_ack_0, ack => convolution3D_CP_3583_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	71 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1384_Update/ca
      -- 
    ca_4087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1384_inst_ack_1, ack => convolution3D_CP_3583_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_Update/cr
      -- 
    ra_4096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1392_inst_ack_0, ack => convolution3D_CP_3583_elements(57)); -- 
    cr_4100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(57), ack => RPIPE_maxpool_input_pipe_1392_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1392_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_Sample/rr
      -- 
    ca_4101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1392_inst_ack_1, ack => convolution3D_CP_3583_elements(58)); -- 
    rr_4109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(58), ack => type_cast_1396_inst_req_0); -- 
    rr_4123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(58), ack => RPIPE_maxpool_input_pipe_1405_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_Sample/ra
      -- 
    ra_4110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1396_inst_ack_0, ack => convolution3D_CP_3583_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	71 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1396_Update/ca
      -- 
    ca_4115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1396_inst_ack_1, ack => convolution3D_CP_3583_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_update_start_
      -- CP-element group 61: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_Update/cr
      -- 
    ra_4124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1405_inst_ack_0, ack => convolution3D_CP_3583_elements(61)); -- 
    cr_4128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(61), ack => RPIPE_maxpool_input_pipe_1405_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/RPIPE_maxpool_input_pipe_1405_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_Sample/rr
      -- 
    ca_4129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1405_inst_ack_1, ack => convolution3D_CP_3583_elements(62)); -- 
    rr_4137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(62), ack => type_cast_1409_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_Sample/ra
      -- 
    ra_4138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1409_inst_ack_0, ack => convolution3D_CP_3583_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	71 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1409_Update/ca
      -- 
    ca_4143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1409_inst_ack_1, ack => convolution3D_CP_3583_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	16 
    -- CP-element group 65: 	12 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_Sample/rr
      -- 
    rr_4151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(65), ack => type_cast_1418_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(16) & convolution3D_CP_3583_elements(12);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_Sample/ra
      -- 
    ra_4152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_0, ack => convolution3D_CP_3583_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1418_Update/ca
      -- 
    ca_4157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_1, ack => convolution3D_CP_3583_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	20 
    -- CP-element group 68: 	24 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_Sample/rr
      -- 
    rr_4165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(68), ack => type_cast_1422_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(20) & convolution3D_CP_3583_elements(24);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_Sample/ra
      -- 
    ra_4166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1422_inst_ack_0, ack => convolution3D_CP_3583_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/type_cast_1422_Update/ca
      -- 
    ca_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1422_inst_ack_1, ack => convolution3D_CP_3583_elements(70)); -- 
    -- CP-element group 71:  branch  join  transition  place  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	52 
    -- CP-element group 71: 	48 
    -- CP-element group 71: 	28 
    -- CP-element group 71: 	40 
    -- CP-element group 71: 	32 
    -- CP-element group 71: 	36 
    -- CP-element group 71: 	44 
    -- CP-element group 71: 	56 
    -- CP-element group 71: 	60 
    -- CP-element group 71: 	64 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: 	4 
    -- CP-element group 71: 	8 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (10) 
      -- CP-element group 71: 	 branch_block_stmt_1215/if_stmt_1440__entry__
      -- CP-element group 71: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439/$exit
      -- CP-element group 71: 	 branch_block_stmt_1215/assign_stmt_1218_to_assign_stmt_1439__exit__
      -- CP-element group 71: 	 branch_block_stmt_1215/if_stmt_1440_dead_link/$entry
      -- CP-element group 71: 	 branch_block_stmt_1215/if_stmt_1440_eval_test/$entry
      -- CP-element group 71: 	 branch_block_stmt_1215/if_stmt_1440_eval_test/$exit
      -- CP-element group 71: 	 branch_block_stmt_1215/if_stmt_1440_eval_test/branch_req
      -- CP-element group 71: 	 branch_block_stmt_1215/R_cmp368_1441_place
      -- CP-element group 71: 	 branch_block_stmt_1215/if_stmt_1440_if_link/$entry
      -- CP-element group 71: 	 branch_block_stmt_1215/if_stmt_1440_else_link/$entry
      -- 
    branch_req_4179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(71), ack => if_stmt_1440_branch_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(52) & convolution3D_CP_3583_elements(48) & convolution3D_CP_3583_elements(28) & convolution3D_CP_3583_elements(40) & convolution3D_CP_3583_elements(32) & convolution3D_CP_3583_elements(36) & convolution3D_CP_3583_elements(44) & convolution3D_CP_3583_elements(56) & convolution3D_CP_3583_elements(60) & convolution3D_CP_3583_elements(64) & convolution3D_CP_3583_elements(67) & convolution3D_CP_3583_elements(70) & convolution3D_CP_3583_elements(4) & convolution3D_CP_3583_elements(8);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: 	75 
    -- CP-element group 72: 	76 
    -- CP-element group 72: 	77 
    -- CP-element group 72: 	80 
    -- CP-element group 72:  members (27) 
      -- CP-element group 72: 	 branch_block_stmt_1215/merge_stmt_1446__exit__
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521__entry__
      -- CP-element group 72: 	 branch_block_stmt_1215/if_stmt_1440_if_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_1215/if_stmt_1440_if_link/if_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_1215/entry_bbx_xnph370
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/$entry
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_update_start_
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_Update/cr
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_update_start_
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_Update/cr
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_update_start_
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_Update/cr
      -- CP-element group 72: 	 branch_block_stmt_1215/entry_bbx_xnph370_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_1215/entry_bbx_xnph370_PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_1215/merge_stmt_1446_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1215/merge_stmt_1446_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_1215/merge_stmt_1446_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_1215/merge_stmt_1446_PhiAck/dummy
      -- 
    if_choice_transition_4184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1440_branch_ack_1, ack => convolution3D_CP_3583_elements(72)); -- 
    rr_4201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(72), ack => type_cast_1471_inst_req_0); -- 
    cr_4206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(72), ack => type_cast_1471_inst_req_1); -- 
    rr_4215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(72), ack => type_cast_1480_inst_req_0); -- 
    cr_4220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(72), ack => type_cast_1480_inst_req_1); -- 
    cr_4234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(72), ack => type_cast_1514_inst_req_1); -- 
    -- CP-element group 73:  transition  place  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	329 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_1215/if_stmt_1440_else_link/$exit
      -- CP-element group 73: 	 branch_block_stmt_1215/if_stmt_1440_else_link/else_choice_transition
      -- CP-element group 73: 	 branch_block_stmt_1215/entry_forx_xend
      -- CP-element group 73: 	 branch_block_stmt_1215/entry_forx_xend_PhiReq/$entry
      -- CP-element group 73: 	 branch_block_stmt_1215/entry_forx_xend_PhiReq/phi_stmt_1707/$entry
      -- CP-element group 73: 	 branch_block_stmt_1215/entry_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/$entry
      -- 
    else_choice_transition_4188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1440_branch_ack_0, ack => convolution3D_CP_3583_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_Sample/ra
      -- 
    ra_4202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1471_inst_ack_0, ack => convolution3D_CP_3583_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	72 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1471_Update/ca
      -- 
    ca_4207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1471_inst_ack_1, ack => convolution3D_CP_3583_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	72 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_Sample/ra
      -- 
    ra_4216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1480_inst_ack_0, ack => convolution3D_CP_3583_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	72 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1480_Update/ca
      -- 
    ca_4221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1480_inst_ack_1, ack => convolution3D_CP_3583_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_Sample/rr
      -- 
    rr_4229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(78), ack => type_cast_1514_inst_req_0); -- 
    convolution3D_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(75) & convolution3D_CP_3583_elements(77);
      gj_convolution3D_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_Sample/ra
      -- 
    ra_4230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1514_inst_ack_0, ack => convolution3D_CP_3583_elements(79)); -- 
    -- CP-element group 80:  transition  place  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	72 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	323 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521__exit__
      -- CP-element group 80: 	 branch_block_stmt_1215/bbx_xnph370_forx_xbody
      -- CP-element group 80: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/$exit
      -- CP-element group 80: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1215/assign_stmt_1451_to_assign_stmt_1521/type_cast_1514_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_1215/bbx_xnph370_forx_xbody_PhiReq/$entry
      -- CP-element group 80: 	 branch_block_stmt_1215/bbx_xnph370_forx_xbody_PhiReq/phi_stmt_1524/$entry
      -- CP-element group 80: 	 branch_block_stmt_1215/bbx_xnph370_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/$entry
      -- 
    ca_4235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1514_inst_ack_1, ack => convolution3D_CP_3583_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	328 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	120 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_final_index_sum_regn_sample_complete
      -- CP-element group 81: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_final_index_sum_regn_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_final_index_sum_regn_Sample/ack
      -- 
    ack_4264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1536_index_offset_ack_0, ack => convolution3D_CP_3583_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	328 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (11) 
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_root_address_calculated
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_offset_calculated
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_final_index_sum_regn_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_final_index_sum_regn_Update/ack
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_base_plus_offset/$entry
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_base_plus_offset/$exit
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_base_plus_offset/sum_rename_req
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_base_plus_offset/sum_rename_ack
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_request/$entry
      -- CP-element group 82: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_request/req
      -- 
    ack_4269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1536_index_offset_ack_1, ack => convolution3D_CP_3583_elements(82)); -- 
    req_4278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(82), ack => addr_of_1537_final_reg_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_request/$exit
      -- CP-element group 83: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_request/ack
      -- 
    ack_4279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1537_final_reg_ack_0, ack => convolution3D_CP_3583_elements(83)); -- 
    -- CP-element group 84:  fork  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	328 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	117 
    -- CP-element group 84:  members (19) 
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_complete/$exit
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_complete/ack
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_base_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_word_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_root_address_calculated
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_base_address_resized
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_base_addr_resize/$entry
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_base_addr_resize/$exit
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_base_addr_resize/base_resize_req
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_base_addr_resize/base_resize_ack
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_base_plus_offset/$entry
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_base_plus_offset/$exit
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_base_plus_offset/sum_rename_req
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_base_plus_offset/sum_rename_ack
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_word_addrgen/$entry
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_word_addrgen/$exit
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_word_addrgen/root_register_req
      -- CP-element group 84: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_word_addrgen/root_register_ack
      -- 
    ack_4284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1537_final_reg_ack_1, ack => convolution3D_CP_3583_elements(84)); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	328 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_update_start_
      -- CP-element group 85: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_Sample/ra
      -- CP-element group 85: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_Update/cr
      -- 
    ra_4293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1540_inst_ack_0, ack => convolution3D_CP_3583_elements(85)); -- 
    cr_4297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(85), ack => RPIPE_maxpool_input_pipe_1540_inst_req_1); -- 
    -- CP-element group 86:  fork  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: 	89 
    -- CP-element group 86:  members (9) 
      -- CP-element group 86: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_Sample/rr
      -- 
    ca_4298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1540_inst_ack_1, ack => convolution3D_CP_3583_elements(86)); -- 
    rr_4306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(86), ack => type_cast_1544_inst_req_0); -- 
    rr_4320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(86), ack => RPIPE_maxpool_input_pipe_1553_inst_req_0); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_Sample/ra
      -- 
    ra_4307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1544_inst_ack_0, ack => convolution3D_CP_3583_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	328 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	117 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_Update/ca
      -- 
    ca_4312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1544_inst_ack_1, ack => convolution3D_CP_3583_elements(88)); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	86 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_update_start_
      -- CP-element group 89: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_Update/cr
      -- 
    ra_4321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1553_inst_ack_0, ack => convolution3D_CP_3583_elements(89)); -- 
    cr_4325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(89), ack => RPIPE_maxpool_input_pipe_1553_inst_req_1); -- 
    -- CP-element group 90:  fork  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: 	93 
    -- CP-element group 90:  members (9) 
      -- CP-element group 90: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1553_Update/ca
      -- CP-element group 90: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_Sample/rr
      -- 
    ca_4326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1553_inst_ack_1, ack => convolution3D_CP_3583_elements(90)); -- 
    rr_4334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(90), ack => type_cast_1557_inst_req_0); -- 
    rr_4348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(90), ack => RPIPE_maxpool_input_pipe_1571_inst_req_0); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_Sample/ra
      -- 
    ra_4335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1557_inst_ack_0, ack => convolution3D_CP_3583_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	328 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	117 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_Update/ca
      -- 
    ca_4340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1557_inst_ack_1, ack => convolution3D_CP_3583_elements(92)); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	90 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_update_start_
      -- CP-element group 93: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_Update/cr
      -- 
    ra_4349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1571_inst_ack_0, ack => convolution3D_CP_3583_elements(93)); -- 
    cr_4353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(93), ack => RPIPE_maxpool_input_pipe_1571_inst_req_1); -- 
    -- CP-element group 94:  fork  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94: 	97 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1571_Update/ca
      -- CP-element group 94: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_Sample/rr
      -- 
    ca_4354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1571_inst_ack_1, ack => convolution3D_CP_3583_elements(94)); -- 
    rr_4376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(94), ack => RPIPE_maxpool_input_pipe_1589_inst_req_0); -- 
    rr_4362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(94), ack => type_cast_1575_inst_req_0); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_Sample/ra
      -- 
    ra_4363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1575_inst_ack_0, ack => convolution3D_CP_3583_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	328 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	117 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_Update/ca
      -- 
    ca_4368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1575_inst_ack_1, ack => convolution3D_CP_3583_elements(96)); -- 
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	94 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_update_start_
      -- CP-element group 97: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_Sample/ra
      -- CP-element group 97: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_Update/cr
      -- 
    ra_4377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1589_inst_ack_0, ack => convolution3D_CP_3583_elements(97)); -- 
    cr_4381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(97), ack => RPIPE_maxpool_input_pipe_1589_inst_req_1); -- 
    -- CP-element group 98:  fork  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	101 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1589_Update/ca
      -- CP-element group 98: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_Sample/rr
      -- 
    ca_4382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1589_inst_ack_1, ack => convolution3D_CP_3583_elements(98)); -- 
    rr_4390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(98), ack => type_cast_1593_inst_req_0); -- 
    rr_4404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(98), ack => RPIPE_maxpool_input_pipe_1607_inst_req_0); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_Sample/ra
      -- 
    ra_4391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1593_inst_ack_0, ack => convolution3D_CP_3583_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	328 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	117 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_Update/ca
      -- 
    ca_4396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1593_inst_ack_1, ack => convolution3D_CP_3583_elements(100)); -- 
    -- CP-element group 101:  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	98 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_update_start_
      -- CP-element group 101: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_Sample/ra
      -- CP-element group 101: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_Update/cr
      -- 
    ra_4405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1607_inst_ack_0, ack => convolution3D_CP_3583_elements(101)); -- 
    cr_4409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(101), ack => RPIPE_maxpool_input_pipe_1607_inst_req_1); -- 
    -- CP-element group 102:  fork  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	105 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (9) 
      -- CP-element group 102: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1607_Update/ca
      -- CP-element group 102: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_Sample/rr
      -- 
    ca_4410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1607_inst_ack_1, ack => convolution3D_CP_3583_elements(102)); -- 
    rr_4432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(102), ack => RPIPE_maxpool_input_pipe_1625_inst_req_0); -- 
    rr_4418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(102), ack => type_cast_1611_inst_req_0); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_Sample/ra
      -- 
    ra_4419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1611_inst_ack_0, ack => convolution3D_CP_3583_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	328 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	117 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_Update/ca
      -- 
    ca_4424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1611_inst_ack_1, ack => convolution3D_CP_3583_elements(104)); -- 
    -- CP-element group 105:  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	102 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (6) 
      -- CP-element group 105: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_update_start_
      -- CP-element group 105: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_Update/cr
      -- 
    ra_4433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1625_inst_ack_0, ack => convolution3D_CP_3583_elements(105)); -- 
    cr_4437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(105), ack => RPIPE_maxpool_input_pipe_1625_inst_req_1); -- 
    -- CP-element group 106:  fork  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106: 	109 
    -- CP-element group 106:  members (9) 
      -- CP-element group 106: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1625_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_Sample/rr
      -- CP-element group 106: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_Sample/rr
      -- 
    ca_4438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1625_inst_ack_1, ack => convolution3D_CP_3583_elements(106)); -- 
    rr_4446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(106), ack => type_cast_1629_inst_req_0); -- 
    rr_4460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(106), ack => RPIPE_maxpool_input_pipe_1643_inst_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_Sample/ra
      -- 
    ra_4447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1629_inst_ack_0, ack => convolution3D_CP_3583_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	328 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	117 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_Update/ca
      -- 
    ca_4452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1629_inst_ack_1, ack => convolution3D_CP_3583_elements(108)); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	106 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_Update/cr
      -- 
    ra_4461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1643_inst_ack_0, ack => convolution3D_CP_3583_elements(109)); -- 
    cr_4465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(109), ack => RPIPE_maxpool_input_pipe_1643_inst_req_1); -- 
    -- CP-element group 110:  fork  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (9) 
      -- CP-element group 110: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1643_Update/ca
      -- CP-element group 110: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_Sample/rr
      -- 
    ca_4466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1643_inst_ack_1, ack => convolution3D_CP_3583_elements(110)); -- 
    rr_4474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(110), ack => type_cast_1647_inst_req_0); -- 
    rr_4488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(110), ack => RPIPE_maxpool_input_pipe_1661_inst_req_0); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_Sample/ra
      -- 
    ra_4475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1647_inst_ack_0, ack => convolution3D_CP_3583_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	328 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	117 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_Update/ca
      -- 
    ca_4480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1647_inst_ack_1, ack => convolution3D_CP_3583_elements(112)); -- 
    -- CP-element group 113:  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (6) 
      -- CP-element group 113: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_update_start_
      -- CP-element group 113: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_Update/cr
      -- 
    ra_4489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1661_inst_ack_0, ack => convolution3D_CP_3583_elements(113)); -- 
    cr_4493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(113), ack => RPIPE_maxpool_input_pipe_1661_inst_req_1); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1661_Update/ca
      -- CP-element group 114: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_Sample/rr
      -- 
    ca_4494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1661_inst_ack_1, ack => convolution3D_CP_3583_elements(114)); -- 
    rr_4502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(114), ack => type_cast_1665_inst_req_0); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_Sample/ra
      -- 
    ra_4503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1665_inst_ack_0, ack => convolution3D_CP_3583_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	328 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_Update/ca
      -- 
    ca_4508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1665_inst_ack_1, ack => convolution3D_CP_3583_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	96 
    -- CP-element group 117: 	104 
    -- CP-element group 117: 	112 
    -- CP-element group 117: 	108 
    -- CP-element group 117: 	100 
    -- CP-element group 117: 	116 
    -- CP-element group 117: 	84 
    -- CP-element group 117: 	88 
    -- CP-element group 117: 	92 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (9) 
      -- CP-element group 117: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/ptr_deref_1673_Split/$entry
      -- CP-element group 117: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/ptr_deref_1673_Split/$exit
      -- CP-element group 117: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/ptr_deref_1673_Split/split_req
      -- CP-element group 117: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/ptr_deref_1673_Split/split_ack
      -- CP-element group 117: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/word_access_start/$entry
      -- CP-element group 117: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/word_access_start/word_0/$entry
      -- CP-element group 117: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/word_access_start/word_0/rr
      -- 
    rr_4546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(117), ack => ptr_deref_1673_store_0_req_0); -- 
    convolution3D_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(96) & convolution3D_CP_3583_elements(104) & convolution3D_CP_3583_elements(112) & convolution3D_CP_3583_elements(108) & convolution3D_CP_3583_elements(100) & convolution3D_CP_3583_elements(116) & convolution3D_CP_3583_elements(84) & convolution3D_CP_3583_elements(88) & convolution3D_CP_3583_elements(92);
      gj_convolution3D_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/word_access_start/$exit
      -- CP-element group 118: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/word_access_start/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Sample/word_access_start/word_0/ra
      -- 
    ra_4547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1673_store_0_ack_0, ack => convolution3D_CP_3583_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	328 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Update/word_access_complete/$exit
      -- CP-element group 119: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Update/word_access_complete/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Update/word_access_complete/word_0/ca
      -- 
    ca_4558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1673_store_0_ack_1, ack => convolution3D_CP_3583_elements(119)); -- 
    -- CP-element group 120:  branch  join  transition  place  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: 	81 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (10) 
      -- CP-element group 120: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686__exit__
      -- CP-element group 120: 	 branch_block_stmt_1215/if_stmt_1687__entry__
      -- CP-element group 120: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/$exit
      -- CP-element group 120: 	 branch_block_stmt_1215/if_stmt_1687_dead_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_1215/if_stmt_1687_eval_test/$entry
      -- CP-element group 120: 	 branch_block_stmt_1215/if_stmt_1687_eval_test/$exit
      -- CP-element group 120: 	 branch_block_stmt_1215/if_stmt_1687_eval_test/branch_req
      -- CP-element group 120: 	 branch_block_stmt_1215/R_exitcond42_1688_place
      -- CP-element group 120: 	 branch_block_stmt_1215/if_stmt_1687_if_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_1215/if_stmt_1687_else_link/$entry
      -- 
    branch_req_4566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(120), ack => if_stmt_1687_branch_req_0); -- 
    convolution3D_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(119) & convolution3D_CP_3583_elements(81);
      gj_convolution3D_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_1215/merge_stmt_1693__exit__
      -- CP-element group 121: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704__entry__
      -- CP-element group 121: 	 branch_block_stmt_1215/if_stmt_1687_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_1215/if_stmt_1687_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_1215/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 121: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/$entry
      -- CP-element group 121: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_update_start_
      -- CP-element group 121: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_1215/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_1215/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_1215/merge_stmt_1693_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_1215/merge_stmt_1693_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_1215/merge_stmt_1693_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_1215/merge_stmt_1693_PhiAck/dummy
      -- 
    if_choice_transition_4571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1687_branch_ack_1, ack => convolution3D_CP_3583_elements(121)); -- 
    rr_4588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(121), ack => type_cast_1703_inst_req_0); -- 
    cr_4593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(121), ack => type_cast_1703_inst_req_1); -- 
    -- CP-element group 122:  fork  transition  place  input  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	324 
    -- CP-element group 122: 	325 
    -- CP-element group 122:  members (12) 
      -- CP-element group 122: 	 branch_block_stmt_1215/if_stmt_1687_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_1215/if_stmt_1687_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_1215/forx_xbody_forx_xbody
      -- CP-element group 122: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/$entry
      -- CP-element group 122: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/$entry
      -- CP-element group 122: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/$entry
      -- CP-element group 122: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/SplitProtocol/$entry
      -- CP-element group 122: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/SplitProtocol/Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/SplitProtocol/Sample/rr
      -- CP-element group 122: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/SplitProtocol/Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1687_branch_ack_0, ack => convolution3D_CP_3583_elements(122)); -- 
    rr_6122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(122), ack => type_cast_1530_inst_req_0); -- 
    cr_6127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(122), ack => type_cast_1530_inst_req_1); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_Sample/ra
      -- 
    ra_4589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1703_inst_ack_0, ack => convolution3D_CP_3583_elements(123)); -- 
    -- CP-element group 124:  fork  transition  place  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	331 
    -- CP-element group 124: 	330 
    -- CP-element group 124:  members (15) 
      -- CP-element group 124: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 124: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704__exit__
      -- CP-element group 124: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/$exit
      -- CP-element group 124: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_1215/assign_stmt_1700_to_assign_stmt_1704/type_cast_1703_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/$entry
      -- CP-element group 124: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/$entry
      -- CP-element group 124: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/$entry
      -- CP-element group 124: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Sample/rr
      -- CP-element group 124: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Update/cr
      -- 
    ca_4594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1703_inst_ack_1, ack => convolution3D_CP_3583_elements(124)); -- 
    rr_6176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(124), ack => type_cast_1710_inst_req_0); -- 
    cr_6181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(124), ack => type_cast_1710_inst_req_1); -- 
    -- CP-element group 125:  transition  place  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	334 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	353 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_1215/forx_xend_ifx_xend
      -- CP-element group 125: 	 branch_block_stmt_1215/if_stmt_1727_if_link/if_choice_transition
      -- CP-element group 125: 	 branch_block_stmt_1215/if_stmt_1727_if_link/$exit
      -- CP-element group 125: 	 branch_block_stmt_1215/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_1215/forx_xend_ifx_xend_PhiReq/$exit
      -- 
    if_choice_transition_4610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1727_branch_ack_1, ack => convolution3D_CP_3583_elements(125)); -- 
    -- CP-element group 126:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	334 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	133 
    -- CP-element group 126: 	135 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126: 	129 
    -- CP-element group 126: 	130 
    -- CP-element group 126:  members (30) 
      -- CP-element group 126: 	 branch_block_stmt_1215/merge_stmt_1733__exit__
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760__entry__
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_update_start_
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_Update/cr
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_update_start_
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_Sample/rr
      -- CP-element group 126: 	 branch_block_stmt_1215/forx_xend_forx_xbodyx_xix_xpreheader
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_Update/cr
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_Sample/rr
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_Update/cr
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_update_start_
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_update_start_
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_Update/cr
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/$entry
      -- CP-element group 126: 	 branch_block_stmt_1215/if_stmt_1727_else_link/else_choice_transition
      -- CP-element group 126: 	 branch_block_stmt_1215/if_stmt_1727_else_link/$exit
      -- CP-element group 126: 	 branch_block_stmt_1215/forx_xend_forx_xbodyx_xix_xpreheader_PhiReq/$entry
      -- CP-element group 126: 	 branch_block_stmt_1215/forx_xend_forx_xbodyx_xix_xpreheader_PhiReq/$exit
      -- CP-element group 126: 	 branch_block_stmt_1215/merge_stmt_1733_PhiReqMerge
      -- CP-element group 126: 	 branch_block_stmt_1215/merge_stmt_1733_PhiAck/$entry
      -- CP-element group 126: 	 branch_block_stmt_1215/merge_stmt_1733_PhiAck/$exit
      -- CP-element group 126: 	 branch_block_stmt_1215/merge_stmt_1733_PhiAck/dummy
      -- 
    else_choice_transition_4614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1727_branch_ack_0, ack => convolution3D_CP_3583_elements(126)); -- 
    cr_4646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(126), ack => type_cast_1745_inst_req_1); -- 
    rr_4641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(126), ack => type_cast_1745_inst_req_0); -- 
    cr_4632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(126), ack => type_cast_1736_inst_req_1); -- 
    rr_4627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(126), ack => type_cast_1736_inst_req_0); -- 
    cr_4674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(126), ack => type_cast_1759_inst_req_1); -- 
    cr_4660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(126), ack => type_cast_1755_inst_req_1); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_Sample/ra
      -- CP-element group 127: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_sample_completed_
      -- 
    ra_4628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1736_inst_ack_0, ack => convolution3D_CP_3583_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	131 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_Update/ca
      -- CP-element group 128: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1736_update_completed_
      -- 
    ca_4633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1736_inst_ack_1, ack => convolution3D_CP_3583_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	126 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_sample_completed_
      -- 
    ra_4642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1745_inst_ack_0, ack => convolution3D_CP_3583_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	126 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1745_update_completed_
      -- 
    ca_4647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1745_inst_ack_1, ack => convolution3D_CP_3583_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	128 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_sample_start_
      -- 
    rr_4655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(131), ack => type_cast_1755_inst_req_0); -- 
    convolution3D_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(128) & convolution3D_CP_3583_elements(130);
      gj_convolution3D_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_Sample/ra
      -- CP-element group 132: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_Sample/$exit
      -- 
    ra_4656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1755_inst_ack_0, ack => convolution3D_CP_3583_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	126 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_Sample/rr
      -- CP-element group 133: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_Update/ca
      -- CP-element group 133: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1755_Update/$exit
      -- 
    ca_4661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1755_inst_ack_1, ack => convolution3D_CP_3583_elements(133)); -- 
    rr_4669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(133), ack => type_cast_1759_inst_req_0); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_Sample/ra
      -- CP-element group 134: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_sample_completed_
      -- 
    ra_4670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1759_inst_ack_0, ack => convolution3D_CP_3583_elements(134)); -- 
    -- CP-element group 135:  fork  transition  place  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	126 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	342 
    -- CP-element group 135: 	343 
    -- CP-element group 135:  members (11) 
      -- CP-element group 135: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760__exit__
      -- CP-element group 135: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi
      -- CP-element group 135: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/type_cast_1759_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_1215/assign_stmt_1737_to_assign_stmt_1760/$exit
      -- CP-element group 135: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 135: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1770/$entry
      -- CP-element group 135: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/$entry
      -- CP-element group 135: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1763/$entry
      -- CP-element group 135: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/$entry
      -- 
    ca_4675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1759_inst_ack_1, ack => convolution3D_CP_3583_elements(135)); -- 
    -- CP-element group 136:  transition  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	348 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (6) 
      -- CP-element group 136: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_Update/cr
      -- CP-element group 136: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_Sample/ra
      -- CP-element group 136: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_update_start_
      -- CP-element group 136: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_sample_completed_
      -- 
    ra_4687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1779_inst_ack_0, ack => convolution3D_CP_3583_elements(136)); -- 
    cr_4691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(136), ack => RPIPE_maxpool_input_pipe_1779_inst_req_1); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_Sample/rr
      -- CP-element group 137: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_Update/ca
      -- CP-element group 137: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_update_completed_
      -- 
    ca_4692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1779_inst_ack_1, ack => convolution3D_CP_3583_elements(137)); -- 
    rr_4700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(137), ack => type_cast_1783_inst_req_0); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_sample_completed_
      -- 
    ra_4701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1783_inst_ack_0, ack => convolution3D_CP_3583_elements(138)); -- 
    -- CP-element group 139:  branch  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	348 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (13) 
      -- CP-element group 139: 	 branch_block_stmt_1215/if_stmt_1807__entry__
      -- CP-element group 139: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806__exit__
      -- CP-element group 139: 	 branch_block_stmt_1215/R_exitcond6_1808_place
      -- CP-element group 139: 	 branch_block_stmt_1215/if_stmt_1807_eval_test/$exit
      -- CP-element group 139: 	 branch_block_stmt_1215/if_stmt_1807_eval_test/$entry
      -- CP-element group 139: 	 branch_block_stmt_1215/if_stmt_1807_dead_link/$entry
      -- CP-element group 139: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_1215/if_stmt_1807_eval_test/branch_req
      -- CP-element group 139: 	 branch_block_stmt_1215/if_stmt_1807_else_link/$entry
      -- CP-element group 139: 	 branch_block_stmt_1215/if_stmt_1807_if_link/$entry
      -- CP-element group 139: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/$exit
      -- 
    ca_4706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1783_inst_ack_1, ack => convolution3D_CP_3583_elements(139)); -- 
    branch_req_4714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(139), ack => if_stmt_1807_branch_req_0); -- 
    -- CP-element group 140:  fork  transition  place  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	349 
    -- CP-element group 140: 	350 
    -- CP-element group 140:  members (12) 
      -- CP-element group 140: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 140: 	 branch_block_stmt_1215/if_stmt_1807_if_link/if_choice_transition
      -- CP-element group 140: 	 branch_block_stmt_1215/if_stmt_1807_if_link/$exit
      -- CP-element group 140: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 140: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/$entry
      -- CP-element group 140: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/$entry
      -- CP-element group 140: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/$entry
      -- CP-element group 140: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/SplitProtocol/$entry
      -- CP-element group 140: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/SplitProtocol/Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/SplitProtocol/Sample/rr
      -- CP-element group 140: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/SplitProtocol/Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1807_branch_ack_1, ack => convolution3D_CP_3583_elements(140)); -- 
    rr_6297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(140), ack => type_cast_1817_inst_req_0); -- 
    cr_6302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(140), ack => type_cast_1817_inst_req_1); -- 
    -- CP-element group 141:  fork  transition  place  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	335 
    -- CP-element group 141: 	336 
    -- CP-element group 141: 	338 
    -- CP-element group 141: 	339 
    -- CP-element group 141:  members (20) 
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 141: 	 branch_block_stmt_1215/if_stmt_1807_else_link/else_choice_transition
      -- CP-element group 141: 	 branch_block_stmt_1215/if_stmt_1807_else_link/$exit
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Sample/rr
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Update/cr
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/SplitProtocol/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/SplitProtocol/Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/SplitProtocol/Sample/rr
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/SplitProtocol/Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1807_branch_ack_0, ack => convolution3D_CP_3583_elements(141)); -- 
    rr_6219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(141), ack => type_cast_1773_inst_req_0); -- 
    cr_6224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(141), ack => type_cast_1773_inst_req_1); -- 
    rr_6242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(141), ack => type_cast_1766_inst_req_0); -- 
    cr_6247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(141), ack => type_cast_1766_inst_req_1); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	352 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_Sample/ra
      -- CP-element group 142: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_sample_completed_
      -- 
    ra_4737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1821_inst_ack_0, ack => convolution3D_CP_3583_elements(142)); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	352 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	148 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_Update/ca
      -- CP-element group 143: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_update_completed_
      -- 
    ca_4742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1821_inst_ack_1, ack => convolution3D_CP_3583_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	352 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	151 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_final_index_sum_regn_Sample/ack
      -- CP-element group 144: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_final_index_sum_regn_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_final_index_sum_regn_sample_complete
      -- 
    ack_4768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1850_index_offset_ack_0, ack => convolution3D_CP_3583_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	352 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (11) 
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_offset_calculated
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_request/req
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_request/$entry
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_base_plus_offset/sum_rename_ack
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_root_address_calculated
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_base_plus_offset/sum_rename_req
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_base_plus_offset/$exit
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_base_plus_offset/$entry
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_final_index_sum_regn_Update/ack
      -- CP-element group 145: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_final_index_sum_regn_Update/$exit
      -- 
    ack_4773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1850_index_offset_ack_1, ack => convolution3D_CP_3583_elements(145)); -- 
    req_4782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(145), ack => addr_of_1851_final_reg_req_0); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_request/$exit
      -- CP-element group 146: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_request/ack
      -- 
    ack_4783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1851_final_reg_ack_0, ack => convolution3D_CP_3583_elements(146)); -- 
    -- CP-element group 147:  fork  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	352 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (19) 
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_base_addr_resize/$entry
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_base_address_resized
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_word_address_calculated
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_root_address_calculated
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_base_address_calculated
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_complete/ack
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_complete/$exit
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_word_addrgen/root_register_ack
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_word_addrgen/root_register_req
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_word_addrgen/$exit
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_word_addrgen/$entry
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_base_plus_offset/sum_rename_ack
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_base_plus_offset/sum_rename_req
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_base_plus_offset/$exit
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_base_plus_offset/$entry
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_base_addr_resize/base_resize_ack
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_base_addr_resize/base_resize_req
      -- CP-element group 147: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_base_addr_resize/$exit
      -- 
    ack_4788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1851_final_reg_ack_1, ack => convolution3D_CP_3583_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: 	143 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148:  members (9) 
      -- CP-element group 148: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/word_access_start/word_0/rr
      -- CP-element group 148: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/word_access_start/word_0/$entry
      -- CP-element group 148: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/ptr_deref_1854_Split/split_req
      -- CP-element group 148: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/ptr_deref_1854_Split/split_ack
      -- CP-element group 148: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/ptr_deref_1854_Split/$exit
      -- CP-element group 148: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/ptr_deref_1854_Split/$entry
      -- CP-element group 148: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/word_access_start/$entry
      -- CP-element group 148: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/$entry
      -- 
    rr_4826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(148), ack => ptr_deref_1854_store_0_req_0); -- 
    convolution3D_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(147) & convolution3D_CP_3583_elements(143);
      gj_convolution3D_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (5) 
      -- CP-element group 149: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/word_access_start/word_0/$exit
      -- CP-element group 149: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/word_access_start/word_0/ra
      -- CP-element group 149: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Sample/word_access_start/$exit
      -- 
    ra_4827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1854_store_0_ack_0, ack => convolution3D_CP_3583_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	352 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (5) 
      -- CP-element group 150: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Update/word_access_complete/$exit
      -- CP-element group 150: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Update/word_access_complete/word_0/ca
      -- CP-element group 150: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Update/word_access_complete/word_0/$exit
      -- 
    ca_4838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1854_store_0_ack_1, ack => convolution3D_CP_3583_elements(150)); -- 
    -- CP-element group 151:  join  transition  place  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: 	144 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	353 
    -- CP-element group 151:  members (5) 
      -- CP-element group 151: 	 branch_block_stmt_1215/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 151: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856__exit__
      -- CP-element group 151: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/$exit
      -- CP-element group 151: 	 branch_block_stmt_1215/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 151: 	 branch_block_stmt_1215/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(150) & convolution3D_CP_3583_elements(144);
      gj_convolution3D_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	353 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_sample_completed_
      -- 
    ra_4850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1861_inst_ack_0, ack => convolution3D_CP_3583_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	353 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	158 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_update_completed_
      -- 
    ca_4855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1861_inst_ack_1, ack => convolution3D_CP_3583_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	353 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_sample_completed_
      -- 
    ra_4864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1865_inst_ack_0, ack => convolution3D_CP_3583_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	353 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	158 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_update_completed_
      -- 
    ca_4869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1865_inst_ack_1, ack => convolution3D_CP_3583_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	353 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_sample_completed_
      -- 
    ra_4878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1869_inst_ack_0, ack => convolution3D_CP_3583_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	353 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_update_completed_
      -- 
    ca_4883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1869_inst_ack_1, ack => convolution3D_CP_3583_elements(157)); -- 
    -- CP-element group 158:  branch  join  transition  place  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	155 
    -- CP-element group 158: 	153 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (10) 
      -- CP-element group 158: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891__exit__
      -- CP-element group 158: 	 branch_block_stmt_1215/if_stmt_1892_dead_link/$entry
      -- CP-element group 158: 	 branch_block_stmt_1215/R_cmp157365_1893_place
      -- CP-element group 158: 	 branch_block_stmt_1215/if_stmt_1892_eval_test/$entry
      -- CP-element group 158: 	 branch_block_stmt_1215/if_stmt_1892__entry__
      -- CP-element group 158: 	 branch_block_stmt_1215/if_stmt_1892_else_link/$entry
      -- CP-element group 158: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/$exit
      -- CP-element group 158: 	 branch_block_stmt_1215/if_stmt_1892_if_link/$entry
      -- CP-element group 158: 	 branch_block_stmt_1215/if_stmt_1892_eval_test/branch_req
      -- CP-element group 158: 	 branch_block_stmt_1215/if_stmt_1892_eval_test/$exit
      -- 
    branch_req_4891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(158), ack => if_stmt_1892_branch_req_0); -- 
    convolution3D_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(155) & convolution3D_CP_3583_elements(153) & convolution3D_CP_3583_elements(157);
      gj_convolution3D_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	163 
    -- CP-element group 159: 	164 
    -- CP-element group 159: 	165 
    -- CP-element group 159: 	171 
    -- CP-element group 159: 	166 
    -- CP-element group 159: 	167 
    -- CP-element group 159: 	168 
    -- CP-element group 159: 	161 
    -- CP-element group 159: 	162 
    -- CP-element group 159:  members (39) 
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_Update/cr
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976__entry__
      -- CP-element group 159: 	 branch_block_stmt_1215/merge_stmt_1898__exit__
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_update_start_
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_update_start_
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/ifx_xend_bbx_xnph
      -- CP-element group 159: 	 branch_block_stmt_1215/if_stmt_1892_if_link/if_choice_transition
      -- CP-element group 159: 	 branch_block_stmt_1215/if_stmt_1892_if_link/$exit
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_Update/cr
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_update_start_
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_Update/cr
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_update_start_
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_Update/cr
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_update_start_
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_Update/cr
      -- CP-element group 159: 	 branch_block_stmt_1215/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 159: 	 branch_block_stmt_1215/merge_stmt_1898_PhiReqMerge
      -- CP-element group 159: 	 branch_block_stmt_1215/merge_stmt_1898_PhiAck/$entry
      -- CP-element group 159: 	 branch_block_stmt_1215/merge_stmt_1898_PhiAck/$exit
      -- CP-element group 159: 	 branch_block_stmt_1215/merge_stmt_1898_PhiAck/dummy
      -- 
    if_choice_transition_4896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1892_branch_ack_1, ack => convolution3D_CP_3583_elements(159)); -- 
    cr_4918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(159), ack => type_cast_1913_inst_req_1); -- 
    rr_4913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(159), ack => type_cast_1913_inst_req_0); -- 
    rr_4927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(159), ack => type_cast_1917_inst_req_0); -- 
    cr_4932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(159), ack => type_cast_1917_inst_req_1); -- 
    rr_4941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(159), ack => type_cast_1926_inst_req_0); -- 
    cr_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(159), ack => type_cast_1926_inst_req_1); -- 
    rr_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(159), ack => type_cast_1935_inst_req_0); -- 
    cr_4960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(159), ack => type_cast_1935_inst_req_1); -- 
    cr_4974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(159), ack => type_cast_1969_inst_req_1); -- 
    -- CP-element group 160:  transition  place  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	363 
    -- CP-element group 160:  members (6) 
      -- CP-element group 160: 	 branch_block_stmt_1215/ifx_xend_forx_xend211
      -- CP-element group 160: 	 branch_block_stmt_1215/if_stmt_1892_else_link/else_choice_transition
      -- CP-element group 160: 	 branch_block_stmt_1215/if_stmt_1892_else_link/$exit
      -- CP-element group 160: 	 branch_block_stmt_1215/ifx_xend_forx_xend211_PhiReq/$entry
      -- CP-element group 160: 	 branch_block_stmt_1215/ifx_xend_forx_xend211_PhiReq/phi_stmt_2162/$entry
      -- CP-element group 160: 	 branch_block_stmt_1215/ifx_xend_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/$entry
      -- 
    else_choice_transition_4900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1892_branch_ack_0, ack => convolution3D_CP_3583_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_Sample/ra
      -- 
    ra_4914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1913_inst_ack_0, ack => convolution3D_CP_3583_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	159 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	169 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_Update/ca
      -- CP-element group 162: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1913_Update/$exit
      -- 
    ca_4919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1913_inst_ack_1, ack => convolution3D_CP_3583_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	159 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_Sample/ra
      -- 
    ra_4928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1917_inst_ack_0, ack => convolution3D_CP_3583_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	159 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	169 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1917_Update/ca
      -- 
    ca_4933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1917_inst_ack_1, ack => convolution3D_CP_3583_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	159 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_Sample/ra
      -- 
    ra_4942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1926_inst_ack_0, ack => convolution3D_CP_3583_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	159 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	169 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1926_Update/ca
      -- 
    ca_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1926_inst_ack_1, ack => convolution3D_CP_3583_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	159 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_Sample/ra
      -- 
    ra_4956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1935_inst_ack_0, ack => convolution3D_CP_3583_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	159 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1935_Update/ca
      -- 
    ca_4961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1935_inst_ack_1, ack => convolution3D_CP_3583_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	164 
    -- CP-element group 169: 	166 
    -- CP-element group 169: 	168 
    -- CP-element group 169: 	162 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_Sample/rr
      -- 
    rr_4969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(169), ack => type_cast_1969_inst_req_0); -- 
    convolution3D_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(164) & convolution3D_CP_3583_elements(166) & convolution3D_CP_3583_elements(168) & convolution3D_CP_3583_elements(162);
      gj_convolution3D_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_Sample/ra
      -- 
    ra_4970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1969_inst_ack_0, ack => convolution3D_CP_3583_elements(170)); -- 
    -- CP-element group 171:  transition  place  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	159 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	354 
    -- CP-element group 171:  members (9) 
      -- CP-element group 171: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/$exit
      -- CP-element group 171: 	 branch_block_stmt_1215/bbx_xnph_forx_xbody159
      -- CP-element group 171: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976__exit__
      -- CP-element group 171: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_1215/assign_stmt_1904_to_assign_stmt_1976/type_cast_1969_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_1215/bbx_xnph_forx_xbody159_PhiReq/$entry
      -- CP-element group 171: 	 branch_block_stmt_1215/bbx_xnph_forx_xbody159_PhiReq/phi_stmt_1979/$entry
      -- CP-element group 171: 	 branch_block_stmt_1215/bbx_xnph_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/$entry
      -- 
    ca_4975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1969_inst_ack_1, ack => convolution3D_CP_3583_elements(171)); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	359 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	211 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_final_index_sum_regn_sample_complete
      -- CP-element group 172: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_final_index_sum_regn_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_final_index_sum_regn_Sample/ack
      -- 
    ack_5004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1991_index_offset_ack_0, ack => convolution3D_CP_3583_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	359 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (11) 
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_root_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_offset_calculated
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_final_index_sum_regn_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_final_index_sum_regn_Update/ack
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_base_plus_offset/$entry
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_base_plus_offset/$exit
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_base_plus_offset/sum_rename_req
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_base_plus_offset/sum_rename_ack
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_request/$entry
      -- CP-element group 173: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_request/req
      -- 
    ack_5009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1991_index_offset_ack_1, ack => convolution3D_CP_3583_elements(173)); -- 
    req_5018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(173), ack => addr_of_1992_final_reg_req_0); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_request/$exit
      -- CP-element group 174: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_request/ack
      -- 
    ack_5019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1992_final_reg_ack_0, ack => convolution3D_CP_3583_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	359 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	208 
    -- CP-element group 175:  members (19) 
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_complete/$exit
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_complete/ack
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_base_address_calculated
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_word_address_calculated
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_root_address_calculated
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_base_address_resized
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_base_addr_resize/$entry
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_base_addr_resize/$exit
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_base_addr_resize/base_resize_req
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_base_addr_resize/base_resize_ack
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_base_plus_offset/$entry
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_base_plus_offset/$exit
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_base_plus_offset/sum_rename_req
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_base_plus_offset/sum_rename_ack
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_word_addrgen/$entry
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_word_addrgen/$exit
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_word_addrgen/root_register_req
      -- CP-element group 175: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_word_addrgen/root_register_ack
      -- 
    ack_5024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1992_final_reg_ack_1, ack => convolution3D_CP_3583_elements(175)); -- 
    -- CP-element group 176:  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	359 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (6) 
      -- CP-element group 176: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_update_start_
      -- CP-element group 176: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_Sample/ra
      -- CP-element group 176: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_Update/cr
      -- 
    ra_5033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1995_inst_ack_0, ack => convolution3D_CP_3583_elements(176)); -- 
    cr_5037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(176), ack => RPIPE_maxpool_input_pipe_1995_inst_req_1); -- 
    -- CP-element group 177:  fork  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: 	180 
    -- CP-element group 177:  members (9) 
      -- CP-element group 177: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_Update/ca
      -- CP-element group 177: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_Sample/rr
      -- CP-element group 177: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_Sample/rr
      -- 
    ca_5038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1995_inst_ack_1, ack => convolution3D_CP_3583_elements(177)); -- 
    rr_5046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(177), ack => type_cast_1999_inst_req_0); -- 
    rr_5060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(177), ack => RPIPE_maxpool_input_pipe_2008_inst_req_0); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_Sample/ra
      -- 
    ra_5047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1999_inst_ack_0, ack => convolution3D_CP_3583_elements(178)); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	359 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	208 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_Update/ca
      -- 
    ca_5052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1999_inst_ack_1, ack => convolution3D_CP_3583_elements(179)); -- 
    -- CP-element group 180:  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	177 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_update_start_
      -- CP-element group 180: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_Sample/ra
      -- CP-element group 180: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_Update/cr
      -- 
    ra_5061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2008_inst_ack_0, ack => convolution3D_CP_3583_elements(180)); -- 
    cr_5065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(180), ack => RPIPE_maxpool_input_pipe_2008_inst_req_1); -- 
    -- CP-element group 181:  fork  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181: 	184 
    -- CP-element group 181:  members (9) 
      -- CP-element group 181: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2008_Update/ca
      -- CP-element group 181: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_Sample/rr
      -- 
    ca_5066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2008_inst_ack_1, ack => convolution3D_CP_3583_elements(181)); -- 
    rr_5074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(181), ack => type_cast_2012_inst_req_0); -- 
    rr_5088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(181), ack => RPIPE_maxpool_input_pipe_2026_inst_req_0); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_Sample/ra
      -- 
    ra_5075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2012_inst_ack_0, ack => convolution3D_CP_3583_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	359 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	208 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_Update/ca
      -- 
    ca_5080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2012_inst_ack_1, ack => convolution3D_CP_3583_elements(183)); -- 
    -- CP-element group 184:  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	181 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (6) 
      -- CP-element group 184: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_Sample/ra
      -- CP-element group 184: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_Update/cr
      -- 
    ra_5089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2026_inst_ack_0, ack => convolution3D_CP_3583_elements(184)); -- 
    cr_5093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(184), ack => RPIPE_maxpool_input_pipe_2026_inst_req_1); -- 
    -- CP-element group 185:  fork  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185: 	188 
    -- CP-element group 185:  members (9) 
      -- CP-element group 185: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2026_Update/ca
      -- CP-element group 185: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_Sample/rr
      -- CP-element group 185: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_Sample/rr
      -- 
    ca_5094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2026_inst_ack_1, ack => convolution3D_CP_3583_elements(185)); -- 
    rr_5102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(185), ack => type_cast_2030_inst_req_0); -- 
    rr_5116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(185), ack => RPIPE_maxpool_input_pipe_2044_inst_req_0); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_Sample/ra
      -- 
    ra_5103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2030_inst_ack_0, ack => convolution3D_CP_3583_elements(186)); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	359 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	208 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_Update/ca
      -- 
    ca_5108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2030_inst_ack_1, ack => convolution3D_CP_3583_elements(187)); -- 
    -- CP-element group 188:  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	185 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (6) 
      -- CP-element group 188: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_update_start_
      -- CP-element group 188: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_Sample/ra
      -- CP-element group 188: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_Update/cr
      -- 
    ra_5117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2044_inst_ack_0, ack => convolution3D_CP_3583_elements(188)); -- 
    cr_5121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(188), ack => RPIPE_maxpool_input_pipe_2044_inst_req_1); -- 
    -- CP-element group 189:  fork  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189: 	192 
    -- CP-element group 189:  members (9) 
      -- CP-element group 189: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2044_Update/ca
      -- CP-element group 189: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_Sample/rr
      -- CP-element group 189: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_Sample/rr
      -- 
    ca_5122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2044_inst_ack_1, ack => convolution3D_CP_3583_elements(189)); -- 
    rr_5130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(189), ack => type_cast_2048_inst_req_0); -- 
    rr_5144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(189), ack => RPIPE_maxpool_input_pipe_2062_inst_req_0); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_Sample/ra
      -- 
    ra_5131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2048_inst_ack_0, ack => convolution3D_CP_3583_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	359 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	208 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_Update/ca
      -- 
    ca_5136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2048_inst_ack_1, ack => convolution3D_CP_3583_elements(191)); -- 
    -- CP-element group 192:  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	189 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (6) 
      -- CP-element group 192: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_update_start_
      -- CP-element group 192: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_Sample/ra
      -- CP-element group 192: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_Update/$entry
      -- CP-element group 192: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_Update/cr
      -- 
    ra_5145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2062_inst_ack_0, ack => convolution3D_CP_3583_elements(192)); -- 
    cr_5149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(192), ack => RPIPE_maxpool_input_pipe_2062_inst_req_1); -- 
    -- CP-element group 193:  fork  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193: 	196 
    -- CP-element group 193:  members (9) 
      -- CP-element group 193: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2062_Update/ca
      -- CP-element group 193: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_Sample/rr
      -- CP-element group 193: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_Sample/rr
      -- 
    ca_5150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2062_inst_ack_1, ack => convolution3D_CP_3583_elements(193)); -- 
    rr_5158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(193), ack => type_cast_2066_inst_req_0); -- 
    rr_5172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(193), ack => RPIPE_maxpool_input_pipe_2080_inst_req_0); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_Sample/ra
      -- 
    ra_5159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2066_inst_ack_0, ack => convolution3D_CP_3583_elements(194)); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	359 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	208 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_Update/ca
      -- 
    ca_5164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2066_inst_ack_1, ack => convolution3D_CP_3583_elements(195)); -- 
    -- CP-element group 196:  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	193 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196:  members (6) 
      -- CP-element group 196: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_update_start_
      -- CP-element group 196: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_Sample/ra
      -- CP-element group 196: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_Update/$entry
      -- CP-element group 196: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_Update/cr
      -- 
    ra_5173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2080_inst_ack_0, ack => convolution3D_CP_3583_elements(196)); -- 
    cr_5177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(196), ack => RPIPE_maxpool_input_pipe_2080_inst_req_1); -- 
    -- CP-element group 197:  fork  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	200 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (9) 
      -- CP-element group 197: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2080_Update/ca
      -- CP-element group 197: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_Sample/rr
      -- CP-element group 197: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_Sample/rr
      -- 
    ca_5178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2080_inst_ack_1, ack => convolution3D_CP_3583_elements(197)); -- 
    rr_5186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(197), ack => type_cast_2084_inst_req_0); -- 
    rr_5200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(197), ack => RPIPE_maxpool_input_pipe_2098_inst_req_0); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_Sample/ra
      -- 
    ra_5187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2084_inst_ack_0, ack => convolution3D_CP_3583_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	359 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	208 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_Update/ca
      -- 
    ca_5192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2084_inst_ack_1, ack => convolution3D_CP_3583_elements(199)); -- 
    -- CP-element group 200:  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	197 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (6) 
      -- CP-element group 200: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_update_start_
      -- CP-element group 200: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_Update/cr
      -- 
    ra_5201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2098_inst_ack_0, ack => convolution3D_CP_3583_elements(200)); -- 
    cr_5205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(200), ack => RPIPE_maxpool_input_pipe_2098_inst_req_1); -- 
    -- CP-element group 201:  fork  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: 	204 
    -- CP-element group 201:  members (9) 
      -- CP-element group 201: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2098_Update/ca
      -- CP-element group 201: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_sample_start_
      -- CP-element group 201: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_Sample/$entry
      -- CP-element group 201: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_Sample/rr
      -- CP-element group 201: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_sample_start_
      -- CP-element group 201: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_Sample/$entry
      -- CP-element group 201: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_Sample/rr
      -- 
    ca_5206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2098_inst_ack_1, ack => convolution3D_CP_3583_elements(201)); -- 
    rr_5214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(201), ack => type_cast_2102_inst_req_0); -- 
    rr_5228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(201), ack => RPIPE_maxpool_input_pipe_2116_inst_req_0); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_sample_completed_
      -- CP-element group 202: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_Sample/ra
      -- 
    ra_5215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2102_inst_ack_0, ack => convolution3D_CP_3583_elements(202)); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	359 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	208 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_Update/ca
      -- 
    ca_5220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2102_inst_ack_1, ack => convolution3D_CP_3583_elements(203)); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	201 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_update_start_
      -- CP-element group 204: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_Sample/ra
      -- CP-element group 204: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_Update/cr
      -- 
    ra_5229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2116_inst_ack_0, ack => convolution3D_CP_3583_elements(204)); -- 
    cr_5233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(204), ack => RPIPE_maxpool_input_pipe_2116_inst_req_1); -- 
    -- CP-element group 205:  transition  input  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (6) 
      -- CP-element group 205: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_2116_Update/ca
      -- CP-element group 205: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_Sample/rr
      -- 
    ca_5234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2116_inst_ack_1, ack => convolution3D_CP_3583_elements(205)); -- 
    rr_5242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(205), ack => type_cast_2120_inst_req_0); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_Sample/ra
      -- 
    ra_5243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2120_inst_ack_0, ack => convolution3D_CP_3583_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	359 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_Update/ca
      -- 
    ca_5248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2120_inst_ack_1, ack => convolution3D_CP_3583_elements(207)); -- 
    -- CP-element group 208:  join  transition  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	187 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	175 
    -- CP-element group 208: 	199 
    -- CP-element group 208: 	179 
    -- CP-element group 208: 	191 
    -- CP-element group 208: 	183 
    -- CP-element group 208: 	195 
    -- CP-element group 208: 	203 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (9) 
      -- CP-element group 208: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/ptr_deref_2128_Split/$entry
      -- CP-element group 208: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/ptr_deref_2128_Split/$exit
      -- CP-element group 208: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/ptr_deref_2128_Split/split_req
      -- CP-element group 208: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/ptr_deref_2128_Split/split_ack
      -- CP-element group 208: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/word_access_start/$entry
      -- CP-element group 208: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/word_access_start/word_0/$entry
      -- CP-element group 208: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/word_access_start/word_0/rr
      -- 
    rr_5286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(208), ack => ptr_deref_2128_store_0_req_0); -- 
    convolution3D_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(187) & convolution3D_CP_3583_elements(207) & convolution3D_CP_3583_elements(175) & convolution3D_CP_3583_elements(199) & convolution3D_CP_3583_elements(179) & convolution3D_CP_3583_elements(191) & convolution3D_CP_3583_elements(183) & convolution3D_CP_3583_elements(195) & convolution3D_CP_3583_elements(203);
      gj_convolution3D_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/word_access_start/$exit
      -- CP-element group 209: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/word_access_start/word_0/$exit
      -- CP-element group 209: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Sample/word_access_start/word_0/ra
      -- 
    ra_5287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2128_store_0_ack_0, ack => convolution3D_CP_3583_elements(209)); -- 
    -- CP-element group 210:  transition  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	359 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (5) 
      -- CP-element group 210: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Update/word_access_complete/$exit
      -- CP-element group 210: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Update/word_access_complete/word_0/$exit
      -- CP-element group 210: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Update/word_access_complete/word_0/ca
      -- 
    ca_5298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2128_store_0_ack_1, ack => convolution3D_CP_3583_elements(210)); -- 
    -- CP-element group 211:  branch  join  transition  place  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	172 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (10) 
      -- CP-element group 211: 	 branch_block_stmt_1215/if_stmt_2142__entry__
      -- CP-element group 211: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141__exit__
      -- CP-element group 211: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/$exit
      -- CP-element group 211: 	 branch_block_stmt_1215/if_stmt_2142_dead_link/$entry
      -- CP-element group 211: 	 branch_block_stmt_1215/if_stmt_2142_eval_test/$entry
      -- CP-element group 211: 	 branch_block_stmt_1215/if_stmt_2142_eval_test/$exit
      -- CP-element group 211: 	 branch_block_stmt_1215/if_stmt_2142_eval_test/branch_req
      -- CP-element group 211: 	 branch_block_stmt_1215/R_exitcond31_2143_place
      -- CP-element group 211: 	 branch_block_stmt_1215/if_stmt_2142_if_link/$entry
      -- CP-element group 211: 	 branch_block_stmt_1215/if_stmt_2142_else_link/$entry
      -- 
    branch_req_5306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(211), ack => if_stmt_2142_branch_req_0); -- 
    convolution3D_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(172) & convolution3D_CP_3583_elements(210);
      gj_convolution3D_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212: 	215 
    -- CP-element group 212:  members (18) 
      -- CP-element group 212: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159__entry__
      -- CP-element group 212: 	 branch_block_stmt_1215/merge_stmt_2148__exit__
      -- CP-element group 212: 	 branch_block_stmt_1215/if_stmt_2142_if_link/$exit
      -- CP-element group 212: 	 branch_block_stmt_1215/if_stmt_2142_if_link/if_choice_transition
      -- CP-element group 212: 	 branch_block_stmt_1215/forx_xbody159_forx_xcond153x_xforx_xend211_crit_edge
      -- CP-element group 212: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/$entry
      -- CP-element group 212: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_update_start_
      -- CP-element group 212: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_Update/cr
      -- CP-element group 212: 	 branch_block_stmt_1215/forx_xbody159_forx_xcond153x_xforx_xend211_crit_edge_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_1215/forx_xbody159_forx_xcond153x_xforx_xend211_crit_edge_PhiReq/$exit
      -- CP-element group 212: 	 branch_block_stmt_1215/merge_stmt_2148_PhiReqMerge
      -- CP-element group 212: 	 branch_block_stmt_1215/merge_stmt_2148_PhiAck/$entry
      -- CP-element group 212: 	 branch_block_stmt_1215/merge_stmt_2148_PhiAck/$exit
      -- CP-element group 212: 	 branch_block_stmt_1215/merge_stmt_2148_PhiAck/dummy
      -- 
    if_choice_transition_5311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2142_branch_ack_1, ack => convolution3D_CP_3583_elements(212)); -- 
    rr_5328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(212), ack => type_cast_2158_inst_req_0); -- 
    cr_5333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(212), ack => type_cast_2158_inst_req_1); -- 
    -- CP-element group 213:  fork  transition  place  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	355 
    -- CP-element group 213: 	356 
    -- CP-element group 213:  members (12) 
      -- CP-element group 213: 	 branch_block_stmt_1215/if_stmt_2142_else_link/$exit
      -- CP-element group 213: 	 branch_block_stmt_1215/if_stmt_2142_else_link/else_choice_transition
      -- CP-element group 213: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159
      -- CP-element group 213: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/$entry
      -- CP-element group 213: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/$entry
      -- CP-element group 213: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/$entry
      -- CP-element group 213: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/$entry
      -- CP-element group 213: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/SplitProtocol/$entry
      -- CP-element group 213: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/SplitProtocol/Sample/$entry
      -- CP-element group 213: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/SplitProtocol/Sample/rr
      -- CP-element group 213: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/SplitProtocol/Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2142_branch_ack_0, ack => convolution3D_CP_3583_elements(213)); -- 
    rr_6362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(213), ack => type_cast_1985_inst_req_0); -- 
    cr_6367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(213), ack => type_cast_1985_inst_req_1); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_sample_completed_
      -- CP-element group 214: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_Sample/ra
      -- 
    ra_5329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2158_inst_ack_0, ack => convolution3D_CP_3583_elements(214)); -- 
    -- CP-element group 215:  fork  transition  place  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	212 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	360 
    -- CP-element group 215: 	361 
    -- CP-element group 215:  members (15) 
      -- CP-element group 215: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211
      -- CP-element group 215: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159__exit__
      -- CP-element group 215: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/$exit
      -- CP-element group 215: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_Update/$exit
      -- CP-element group 215: 	 branch_block_stmt_1215/assign_stmt_2155_to_assign_stmt_2159/type_cast_2158_Update/ca
      -- CP-element group 215: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/$entry
      -- CP-element group 215: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/$entry
      -- CP-element group 215: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/$entry
      -- CP-element group 215: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/$entry
      -- CP-element group 215: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/SplitProtocol/$entry
      -- CP-element group 215: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/SplitProtocol/Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/SplitProtocol/Sample/rr
      -- CP-element group 215: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/SplitProtocol/Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/SplitProtocol/Update/cr
      -- 
    ca_5334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2158_inst_ack_1, ack => convolution3D_CP_3583_elements(215)); -- 
    rr_6405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(215), ack => type_cast_2165_inst_req_0); -- 
    cr_6410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(215), ack => type_cast_2165_inst_req_1); -- 
    -- CP-element group 216:  transition  place  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	365 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	384 
    -- CP-element group 216:  members (5) 
      -- CP-element group 216: 	 branch_block_stmt_1215/if_stmt_2182_if_link/$exit
      -- CP-element group 216: 	 branch_block_stmt_1215/if_stmt_2182_if_link/if_choice_transition
      -- CP-element group 216: 	 branch_block_stmt_1215/forx_xend211_ifx_xend223
      -- CP-element group 216: 	 branch_block_stmt_1215/forx_xend211_ifx_xend223_PhiReq/$entry
      -- CP-element group 216: 	 branch_block_stmt_1215/forx_xend211_ifx_xend223_PhiReq/$exit
      -- 
    if_choice_transition_5350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2182_branch_ack_1, ack => convolution3D_CP_3583_elements(216)); -- 
    -- CP-element group 217:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	365 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: 	221 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (21) 
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211__entry__
      -- CP-element group 217: 	 branch_block_stmt_1215/merge_stmt_2188__exit__
      -- CP-element group 217: 	 branch_block_stmt_1215/if_stmt_2182_else_link/$exit
      -- CP-element group 217: 	 branch_block_stmt_1215/if_stmt_2182_else_link/else_choice_transition
      -- CP-element group 217: 	 branch_block_stmt_1215/forx_xend211_forx_xbodyx_xi356x_xpreheader
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/$entry
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_sample_start_
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_update_start_
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_Sample/$entry
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_Sample/rr
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_Update/cr
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_update_start_
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_Update/cr
      -- CP-element group 217: 	 branch_block_stmt_1215/forx_xend211_forx_xbodyx_xi356x_xpreheader_PhiReq/$entry
      -- CP-element group 217: 	 branch_block_stmt_1215/forx_xend211_forx_xbodyx_xi356x_xpreheader_PhiReq/$exit
      -- CP-element group 217: 	 branch_block_stmt_1215/merge_stmt_2188_PhiReqMerge
      -- CP-element group 217: 	 branch_block_stmt_1215/merge_stmt_2188_PhiAck/$entry
      -- CP-element group 217: 	 branch_block_stmt_1215/merge_stmt_2188_PhiAck/$exit
      -- CP-element group 217: 	 branch_block_stmt_1215/merge_stmt_2188_PhiAck/dummy
      -- 
    else_choice_transition_5354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2182_branch_ack_0, ack => convolution3D_CP_3583_elements(217)); -- 
    rr_5367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(217), ack => type_cast_2206_inst_req_0); -- 
    cr_5372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(217), ack => type_cast_2206_inst_req_1); -- 
    cr_5386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(217), ack => type_cast_2210_inst_req_1); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_sample_completed_
      -- CP-element group 218: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_Sample/$exit
      -- CP-element group 218: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_Sample/ra
      -- 
    ra_5368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2206_inst_ack_0, ack => convolution3D_CP_3583_elements(218)); -- 
    -- CP-element group 219:  transition  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (6) 
      -- CP-element group 219: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_update_completed_
      -- CP-element group 219: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_Update/$exit
      -- CP-element group 219: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2206_Update/ca
      -- CP-element group 219: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_Sample/rr
      -- 
    ca_5373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2206_inst_ack_1, ack => convolution3D_CP_3583_elements(219)); -- 
    rr_5381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(219), ack => type_cast_2210_inst_req_0); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_Sample/ra
      -- 
    ra_5382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2210_inst_ack_0, ack => convolution3D_CP_3583_elements(220)); -- 
    -- CP-element group 221:  fork  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	217 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	373 
    -- CP-element group 221: 	374 
    -- CP-element group 221:  members (11) 
      -- CP-element group 221: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211__exit__
      -- CP-element group 221: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356
      -- CP-element group 221: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/$exit
      -- CP-element group 221: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_1215/assign_stmt_2193_to_assign_stmt_2211/type_cast_2210_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/$entry
      -- CP-element group 221: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/$entry
      -- CP-element group 221: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/$entry
      -- CP-element group 221: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/$entry
      -- 
    ca_5387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2210_inst_ack_1, ack => convolution3D_CP_3583_elements(221)); -- 
    -- CP-element group 222:  transition  input  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	379 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (6) 
      -- CP-element group 222: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_sample_completed_
      -- CP-element group 222: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_update_start_
      -- CP-element group 222: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_Sample/ra
      -- CP-element group 222: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_Update/$entry
      -- CP-element group 222: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_Update/cr
      -- 
    ra_5399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2230_inst_ack_0, ack => convolution3D_CP_3583_elements(222)); -- 
    cr_5403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(222), ack => RPIPE_maxpool_input_pipe_2230_inst_req_1); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (6) 
      -- CP-element group 223: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_update_completed_
      -- CP-element group 223: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_Update/ca
      -- CP-element group 223: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_Sample/$entry
      -- CP-element group 223: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_Sample/rr
      -- 
    ca_5404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2230_inst_ack_1, ack => convolution3D_CP_3583_elements(223)); -- 
    rr_5412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(223), ack => type_cast_2234_inst_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_Sample/ra
      -- 
    ra_5413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2234_inst_ack_0, ack => convolution3D_CP_3583_elements(224)); -- 
    -- CP-element group 225:  branch  transition  place  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	379 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (13) 
      -- CP-element group 225: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257__exit__
      -- CP-element group 225: 	 branch_block_stmt_1215/if_stmt_2258__entry__
      -- CP-element group 225: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/$exit
      -- CP-element group 225: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_Update/ca
      -- CP-element group 225: 	 branch_block_stmt_1215/if_stmt_2258_dead_link/$entry
      -- CP-element group 225: 	 branch_block_stmt_1215/if_stmt_2258_eval_test/$entry
      -- CP-element group 225: 	 branch_block_stmt_1215/if_stmt_2258_eval_test/$exit
      -- CP-element group 225: 	 branch_block_stmt_1215/if_stmt_2258_eval_test/branch_req
      -- CP-element group 225: 	 branch_block_stmt_1215/R_exitcond_2259_place
      -- CP-element group 225: 	 branch_block_stmt_1215/if_stmt_2258_if_link/$entry
      -- CP-element group 225: 	 branch_block_stmt_1215/if_stmt_2258_else_link/$entry
      -- 
    ca_5418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2234_inst_ack_1, ack => convolution3D_CP_3583_elements(225)); -- 
    branch_req_5426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(225), ack => if_stmt_2258_branch_req_0); -- 
    -- CP-element group 226:  fork  transition  place  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	380 
    -- CP-element group 226: 	381 
    -- CP-element group 226:  members (12) 
      -- CP-element group 226: 	 branch_block_stmt_1215/if_stmt_2258_if_link/$exit
      -- CP-element group 226: 	 branch_block_stmt_1215/if_stmt_2258_if_link/if_choice_transition
      -- CP-element group 226: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363
      -- CP-element group 226: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/$entry
      -- CP-element group 226: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/$entry
      -- CP-element group 226: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/$entry
      -- CP-element group 226: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/$entry
      -- CP-element group 226: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/SplitProtocol/$entry
      -- CP-element group 226: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/SplitProtocol/Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/SplitProtocol/Sample/rr
      -- CP-element group 226: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/SplitProtocol/Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2258_branch_ack_1, ack => convolution3D_CP_3583_elements(226)); -- 
    rr_6537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(226), ack => type_cast_2268_inst_req_0); -- 
    cr_6542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(226), ack => type_cast_2268_inst_req_1); -- 
    -- CP-element group 227:  fork  transition  place  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	366 
    -- CP-element group 227: 	367 
    -- CP-element group 227: 	369 
    -- CP-element group 227: 	370 
    -- CP-element group 227:  members (20) 
      -- CP-element group 227: 	 branch_block_stmt_1215/if_stmt_2258_else_link/$exit
      -- CP-element group 227: 	 branch_block_stmt_1215/if_stmt_2258_else_link/else_choice_transition
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/SplitProtocol/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/SplitProtocol/Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/SplitProtocol/Sample/rr
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/SplitProtocol/Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/SplitProtocol/Update/cr
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/SplitProtocol/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/SplitProtocol/Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/SplitProtocol/Sample/rr
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/SplitProtocol/Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2258_branch_ack_0, ack => convolution3D_CP_3583_elements(227)); -- 
    rr_6459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(227), ack => type_cast_2227_inst_req_0); -- 
    cr_6464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(227), ack => type_cast_2227_inst_req_1); -- 
    rr_6482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(227), ack => type_cast_2220_inst_req_0); -- 
    cr_6487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(227), ack => type_cast_2220_inst_req_1); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	383 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_Sample/ra
      -- CP-element group 228: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_sample_completed_
      -- 
    ra_5449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2272_inst_ack_0, ack => convolution3D_CP_3583_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	383 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	234 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_Update/ca
      -- CP-element group 229: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_update_completed_
      -- 
    ca_5454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2272_inst_ack_1, ack => convolution3D_CP_3583_elements(229)); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	383 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	237 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_final_index_sum_regn_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_final_index_sum_regn_Sample/ack
      -- CP-element group 230: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_final_index_sum_regn_sample_complete
      -- 
    ack_5480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2301_index_offset_ack_0, ack => convolution3D_CP_3583_elements(230)); -- 
    -- CP-element group 231:  transition  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	383 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (11) 
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_offset_calculated
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_root_address_calculated
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_final_index_sum_regn_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_request/req
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_request/$entry
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_base_plus_offset/sum_rename_ack
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_base_plus_offset/sum_rename_req
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_base_plus_offset/$exit
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_base_plus_offset/$entry
      -- CP-element group 231: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_final_index_sum_regn_Update/ack
      -- 
    ack_5485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2301_index_offset_ack_1, ack => convolution3D_CP_3583_elements(231)); -- 
    req_5494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(231), ack => addr_of_2302_final_reg_req_0); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_request/ack
      -- CP-element group 232: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_request/$exit
      -- 
    ack_5495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2302_final_reg_ack_0, ack => convolution3D_CP_3583_elements(232)); -- 
    -- CP-element group 233:  fork  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	383 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (19) 
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_complete/ack
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_base_address_calculated
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_word_address_calculated
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_root_address_calculated
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_base_address_resized
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_base_addr_resize/$entry
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_base_addr_resize/$exit
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_base_addr_resize/base_resize_req
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_base_addr_resize/base_resize_ack
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_base_plus_offset/$entry
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_base_plus_offset/$exit
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_base_plus_offset/sum_rename_req
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_base_plus_offset/sum_rename_ack
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_word_addrgen/$entry
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_complete/$exit
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_word_addrgen/root_register_ack
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_word_addrgen/root_register_req
      -- CP-element group 233: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_word_addrgen/$exit
      -- 
    ack_5500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2302_final_reg_ack_1, ack => convolution3D_CP_3583_elements(233)); -- 
    -- CP-element group 234:  join  transition  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: 	229 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (9) 
      -- CP-element group 234: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/ptr_deref_2305_Split/$entry
      -- CP-element group 234: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/ptr_deref_2305_Split/$exit
      -- CP-element group 234: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/word_access_start/word_0/rr
      -- CP-element group 234: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/word_access_start/word_0/$entry
      -- CP-element group 234: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/word_access_start/$entry
      -- CP-element group 234: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/ptr_deref_2305_Split/split_ack
      -- CP-element group 234: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/ptr_deref_2305_Split/split_req
      -- 
    rr_5538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(234), ack => ptr_deref_2305_store_0_req_0); -- 
    convolution3D_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(233) & convolution3D_CP_3583_elements(229);
      gj_convolution3D_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235:  members (5) 
      -- CP-element group 235: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/word_access_start/word_0/ra
      -- CP-element group 235: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/word_access_start/word_0/$exit
      -- CP-element group 235: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Sample/word_access_start/$exit
      -- 
    ra_5539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2305_store_0_ack_0, ack => convolution3D_CP_3583_elements(235)); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	383 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (5) 
      -- CP-element group 236: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Update/word_access_complete/word_0/ca
      -- CP-element group 236: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Update/word_access_complete/word_0/$exit
      -- CP-element group 236: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Update/word_access_complete/$exit
      -- CP-element group 236: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Update/$exit
      -- 
    ca_5550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2305_store_0_ack_1, ack => convolution3D_CP_3583_elements(236)); -- 
    -- CP-element group 237:  join  transition  place  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: 	230 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	384 
    -- CP-element group 237:  members (5) 
      -- CP-element group 237: 	 branch_block_stmt_1215/getRemainingElementsx_xexit363_ifx_xend223
      -- CP-element group 237: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307__exit__
      -- CP-element group 237: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/$exit
      -- CP-element group 237: 	 branch_block_stmt_1215/getRemainingElementsx_xexit363_ifx_xend223_PhiReq/$entry
      -- CP-element group 237: 	 branch_block_stmt_1215/getRemainingElementsx_xexit363_ifx_xend223_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(236) & convolution3D_CP_3583_elements(230);
      gj_convolution3D_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	384 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_Sample/cra
      -- CP-element group 238: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_sample_completed_
      -- 
    cra_5562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2312_call_ack_0, ack => convolution3D_CP_3583_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	384 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	246 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_Update/cca
      -- CP-element group 239: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_update_completed_
      -- 
    cca_5567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2312_call_ack_1, ack => convolution3D_CP_3583_elements(239)); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	384 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_Update/req
      -- CP-element group 240: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_Update/$entry
      -- CP-element group 240: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_Sample/ack
      -- CP-element group 240: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_update_start_
      -- CP-element group 240: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_sample_completed_
      -- 
    ack_5576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2313_inst_ack_0, ack => convolution3D_CP_3583_elements(240)); -- 
    req_5580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(240), ack => WPIPE_output_pipe_2313_inst_req_1); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_Update/ack
      -- CP-element group 241: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_Sample/req
      -- CP-element group 241: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_update_completed_
      -- 
    ack_5581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2313_inst_ack_1, ack => convolution3D_CP_3583_elements(241)); -- 
    req_5589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(241), ack => WPIPE_output_pipe_2316_inst_req_0); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_sample_completed_
      -- CP-element group 242: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_update_start_
      -- CP-element group 242: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_Sample/ack
      -- CP-element group 242: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_Update/req
      -- 
    ack_5590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2316_inst_ack_0, ack => convolution3D_CP_3583_elements(242)); -- 
    req_5594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(242), ack => WPIPE_output_pipe_2316_inst_req_1); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2316_Update/ack
      -- CP-element group 243: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_Sample/req
      -- 
    ack_5595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2316_inst_ack_1, ack => convolution3D_CP_3583_elements(243)); -- 
    req_5603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(243), ack => WPIPE_output_pipe_2319_inst_req_0); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_update_start_
      -- CP-element group 244: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_Sample/ack
      -- CP-element group 244: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_Update/req
      -- 
    ack_5604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2319_inst_ack_0, ack => convolution3D_CP_3583_elements(244)); -- 
    req_5608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(244), ack => WPIPE_output_pipe_2319_inst_req_1); -- 
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2319_Update/ack
      -- 
    ack_5609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2319_inst_ack_1, ack => convolution3D_CP_3583_elements(245)); -- 
    -- CP-element group 246:  join  fork  transition  place  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	239 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	252 
    -- CP-element group 246: 	247 
    -- CP-element group 246: 	248 
    -- CP-element group 246: 	249 
    -- CP-element group 246: 	250 
    -- CP-element group 246: 	251 
    -- CP-element group 246:  members (22) 
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356__entry__
      -- CP-element group 246: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321__exit__
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_Update/cr
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_Sample/rr
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_update_start_
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_Update/cr
      -- CP-element group 246: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/$exit
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_Sample/rr
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_update_start_
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_Update/cr
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_update_start_
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_Sample/rr
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/$entry
      -- CP-element group 246: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_Sample/$entry
      -- 
    cr_5653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(246), ack => type_cast_2350_inst_req_1); -- 
    rr_5648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(246), ack => type_cast_2350_inst_req_0); -- 
    cr_5639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(246), ack => type_cast_2341_inst_req_1); -- 
    rr_5634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(246), ack => type_cast_2341_inst_req_0); -- 
    cr_5625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(246), ack => type_cast_2331_inst_req_1); -- 
    rr_5620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(246), ack => type_cast_2331_inst_req_0); -- 
    convolution3D_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(239) & convolution3D_CP_3583_elements(245);
      gj_convolution3D_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_Sample/ra
      -- CP-element group 247: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_Sample/$exit
      -- 
    ra_5621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2331_inst_ack_0, ack => convolution3D_CP_3583_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	253 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_Update/ca
      -- CP-element group 248: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2331_update_completed_
      -- 
    ca_5626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2331_inst_ack_1, ack => convolution3D_CP_3583_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	246 
    -- CP-element group 249: successors 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_Sample/ra
      -- CP-element group 249: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_sample_completed_
      -- 
    ra_5635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_0, ack => convolution3D_CP_3583_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	246 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	253 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_Update/ca
      -- CP-element group 250: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2341_update_completed_
      -- 
    ca_5640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_1, ack => convolution3D_CP_3583_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	246 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_Sample/ra
      -- CP-element group 251: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_sample_completed_
      -- 
    ra_5649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2350_inst_ack_0, ack => convolution3D_CP_3583_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	246 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_Update/ca
      -- CP-element group 252: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/type_cast_2350_update_completed_
      -- 
    ca_5654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2350_inst_ack_1, ack => convolution3D_CP_3583_elements(252)); -- 
    -- CP-element group 253:  join  transition  place  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: 	248 
    -- CP-element group 253: 	250 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	385 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356__exit__
      -- CP-element group 253: 	 branch_block_stmt_1215/ifx_xend223_whilex_xbody
      -- CP-element group 253: 	 branch_block_stmt_1215/assign_stmt_2328_to_assign_stmt_2356/$exit
      -- CP-element group 253: 	 branch_block_stmt_1215/ifx_xend223_whilex_xbody_PhiReq/$entry
      -- CP-element group 253: 	 branch_block_stmt_1215/ifx_xend223_whilex_xbody_PhiReq/phi_stmt_2359/$entry
      -- CP-element group 253: 	 branch_block_stmt_1215/ifx_xend223_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/$entry
      -- 
    convolution3D_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(252) & convolution3D_CP_3583_elements(248) & convolution3D_CP_3583_elements(250);
      gj_convolution3D_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	390 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_Update/req
      -- CP-element group 254: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_Sample/ack
      -- CP-element group 254: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_update_start_
      -- CP-element group 254: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_sample_completed_
      -- 
    ack_5666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2372_inst_ack_0, ack => convolution3D_CP_3583_elements(254)); -- 
    req_5670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(254), ack => WPIPE_num_out_pipe_2372_inst_req_1); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_Update/ack
      -- CP-element group 255: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_sample_start_
      -- CP-element group 255: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_Sample/req
      -- CP-element group 255: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_update_completed_
      -- 
    ack_5671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2372_inst_ack_1, ack => convolution3D_CP_3583_elements(255)); -- 
    req_5679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(255), ack => WPIPE_num_out_pipe_2375_inst_req_0); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_update_start_
      -- CP-element group 256: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_Update/req
      -- CP-element group 256: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_Sample/ack
      -- 
    ack_5680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2375_inst_ack_0, ack => convolution3D_CP_3583_elements(256)); -- 
    req_5684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(256), ack => WPIPE_num_out_pipe_2375_inst_req_1); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	262 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_Update/ack
      -- CP-element group 257: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2375_Update/$exit
      -- 
    ack_5685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2375_inst_ack_1, ack => convolution3D_CP_3583_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	390 
    -- CP-element group 258: successors 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_Sample/cra
      -- CP-element group 258: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_sample_completed_
      -- 
    cra_5694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2386_call_ack_0, ack => convolution3D_CP_3583_elements(258)); -- 
    -- CP-element group 259:  transition  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	390 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	262 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_Update/cca
      -- CP-element group 259: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_update_completed_
      -- 
    cca_5699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2386_call_ack_1, ack => convolution3D_CP_3583_elements(259)); -- 
    -- CP-element group 260:  transition  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	390 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_Sample/cra
      -- CP-element group 260: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_sample_completed_
      -- 
    cra_5708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2390_call_ack_0, ack => convolution3D_CP_3583_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	390 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_Update/cca
      -- CP-element group 261: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_update_completed_
      -- 
    cca_5713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2390_call_ack_1, ack => convolution3D_CP_3583_elements(261)); -- 
    -- CP-element group 262:  branch  join  transition  place  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	257 
    -- CP-element group 262: 	259 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (10) 
      -- CP-element group 262: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401__exit__
      -- CP-element group 262: 	 branch_block_stmt_1215/if_stmt_2402__entry__
      -- CP-element group 262: 	 branch_block_stmt_1215/if_stmt_2402_eval_test/$entry
      -- CP-element group 262: 	 branch_block_stmt_1215/if_stmt_2402_eval_test/$exit
      -- CP-element group 262: 	 branch_block_stmt_1215/if_stmt_2402_eval_test/branch_req
      -- CP-element group 262: 	 branch_block_stmt_1215/if_stmt_2402_if_link/$entry
      -- CP-element group 262: 	 branch_block_stmt_1215/if_stmt_2402_else_link/$entry
      -- CP-element group 262: 	 branch_block_stmt_1215/if_stmt_2402_dead_link/$entry
      -- CP-element group 262: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/$exit
      -- CP-element group 262: 	 branch_block_stmt_1215/R_exitcond12_2403_place
      -- 
    branch_req_5721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(262), ack => if_stmt_2402_branch_req_0); -- 
    convolution3D_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(257) & convolution3D_CP_3583_elements(259) & convolution3D_CP_3583_elements(261);
      gj_convolution3D_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	265 
    -- CP-element group 263: 	266 
    -- CP-element group 263: 	267 
    -- CP-element group 263:  members (21) 
      -- CP-element group 263: 	 branch_block_stmt_1215/merge_stmt_2408__exit__
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417__entry__
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_1215/if_stmt_2402_if_link/$exit
      -- CP-element group 263: 	 branch_block_stmt_1215/if_stmt_2402_if_link/if_choice_transition
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_Sample/rr
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_update_start_
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/$entry
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_Update/cr
      -- CP-element group 263: 	 branch_block_stmt_1215/whilex_xbody_whilex_xend
      -- CP-element group 263: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_Sample/rr
      -- CP-element group 263: 	 branch_block_stmt_1215/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 263: 	 branch_block_stmt_1215/merge_stmt_2408_PhiAck/dummy
      -- CP-element group 263: 	 branch_block_stmt_1215/merge_stmt_2408_PhiAck/$exit
      -- CP-element group 263: 	 branch_block_stmt_1215/merge_stmt_2408_PhiAck/$entry
      -- CP-element group 263: 	 branch_block_stmt_1215/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 263: 	 branch_block_stmt_1215/merge_stmt_2408_PhiReqMerge
      -- 
    if_choice_transition_5726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2402_branch_ack_1, ack => convolution3D_CP_3583_elements(263)); -- 
    rr_5743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(263), ack => type_cast_2413_inst_req_0); -- 
    cr_5748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(263), ack => type_cast_2413_inst_req_1); -- 
    rr_5757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(263), ack => RPIPE_input_done_pipe_2416_inst_req_0); -- 
    -- CP-element group 264:  fork  transition  place  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	387 
    -- CP-element group 264: 	386 
    -- CP-element group 264:  members (12) 
      -- CP-element group 264: 	 branch_block_stmt_1215/if_stmt_2402_else_link/else_choice_transition
      -- CP-element group 264: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody
      -- CP-element group 264: 	 branch_block_stmt_1215/if_stmt_2402_else_link/$exit
      -- CP-element group 264: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 264: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/$entry
      -- CP-element group 264: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/$entry
      -- CP-element group 264: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/$entry
      -- CP-element group 264: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/SplitProtocol/$entry
      -- CP-element group 264: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/SplitProtocol/Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/SplitProtocol/Sample/rr
      -- CP-element group 264: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/SplitProtocol/Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2402_branch_ack_0, ack => convolution3D_CP_3583_elements(264)); -- 
    rr_6590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(264), ack => type_cast_2365_inst_req_0); -- 
    cr_6595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(264), ack => type_cast_2365_inst_req_1); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_Sample/ra
      -- CP-element group 265: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_sample_completed_
      -- 
    ra_5744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2413_inst_ack_0, ack => convolution3D_CP_3583_elements(265)); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	263 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	269 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/type_cast_2413_Update/ca
      -- 
    ca_5749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2413_inst_ack_1, ack => convolution3D_CP_3583_elements(266)); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	263 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_update_start_
      -- CP-element group 267: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_Update/cr
      -- CP-element group 267: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_Sample/ra
      -- 
    ra_5758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2416_inst_ack_0, ack => convolution3D_CP_3583_elements(267)); -- 
    cr_5762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(267), ack => RPIPE_input_done_pipe_2416_inst_req_1); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_Update/ca
      -- CP-element group 268: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/RPIPE_input_done_pipe_2416_Update/$exit
      -- 
    ca_5763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2416_inst_ack_1, ack => convolution3D_CP_3583_elements(268)); -- 
    -- CP-element group 269:  join  transition  place  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: 	266 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (7) 
      -- CP-element group 269: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417__exit__
      -- CP-element group 269: 	 branch_block_stmt_1215/assign_stmt_2421__entry__
      -- CP-element group 269: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_Sample/rr
      -- CP-element group 269: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_1215/assign_stmt_2414_to_assign_stmt_2417/$exit
      -- CP-element group 269: 	 branch_block_stmt_1215/assign_stmt_2421/$entry
      -- 
    rr_5774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(269), ack => RPIPE_input_done_pipe_2420_inst_req_0); -- 
    convolution3D_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(268) & convolution3D_CP_3583_elements(266);
      gj_convolution3D_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_Update/cr
      -- CP-element group 270: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_Sample/ra
      -- CP-element group 270: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_update_start_
      -- CP-element group 270: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_sample_completed_
      -- 
    ra_5775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2420_inst_ack_0, ack => convolution3D_CP_3583_elements(270)); -- 
    cr_5779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(270), ack => RPIPE_input_done_pipe_2420_inst_req_1); -- 
    -- CP-element group 271:  fork  transition  place  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	282 
    -- CP-element group 271: 	278 
    -- CP-element group 271: 	279 
    -- CP-element group 271: 	272 
    -- CP-element group 271: 	273 
    -- CP-element group 271: 	275 
    -- CP-element group 271: 	276 
    -- CP-element group 271: 	277 
    -- CP-element group 271:  members (31) 
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454__entry__
      -- CP-element group 271: 	 branch_block_stmt_1215/assign_stmt_2421__exit__
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_update_start_
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_Sample/crr
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_Sample/rr
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/$entry
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_update_start_
      -- CP-element group 271: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_Update/ca
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_Update/ccr
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_Sample/rr
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_update_start_
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_1215/assign_stmt_2421/RPIPE_input_done_pipe_2420_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_update_start_
      -- CP-element group 271: 	 branch_block_stmt_1215/assign_stmt_2421/$exit
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_update_start_
      -- CP-element group 271: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_Update/ccr
      -- 
    ca_5780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2420_inst_ack_1, ack => convolution3D_CP_3583_elements(271)); -- 
    cr_5838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(271), ack => type_cast_2441_inst_req_1); -- 
    crr_5791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(271), ack => call_stmt_2424_call_req_0); -- 
    rr_5833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(271), ack => type_cast_2441_inst_req_0); -- 
    cr_5824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(271), ack => type_cast_2437_inst_req_1); -- 
    ccr_5852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(271), ack => call_stmt_2454_call_req_1); -- 
    rr_5819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(271), ack => type_cast_2437_inst_req_0); -- 
    cr_5810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(271), ack => type_cast_2428_inst_req_1); -- 
    ccr_5796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(271), ack => call_stmt_2424_call_req_1); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_Sample/cra
      -- 
    cra_5792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2424_call_ack_0, ack => convolution3D_CP_3583_elements(272)); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_Sample/rr
      -- CP-element group 273: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_sample_start_
      -- CP-element group 273: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2424_Update/cca
      -- 
    cca_5797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2424_call_ack_1, ack => convolution3D_CP_3583_elements(273)); -- 
    rr_5805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(273), ack => type_cast_2428_inst_req_0); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_Sample/ra
      -- CP-element group 274: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_sample_completed_
      -- 
    ra_5806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2428_inst_ack_0, ack => convolution3D_CP_3583_elements(274)); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	271 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	283 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_Update/ca
      -- CP-element group 275: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2428_update_completed_
      -- 
    ca_5811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2428_inst_ack_1, ack => convolution3D_CP_3583_elements(275)); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	271 
    -- CP-element group 276: successors 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_Sample/ra
      -- CP-element group 276: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_sample_completed_
      -- 
    ra_5820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2437_inst_ack_0, ack => convolution3D_CP_3583_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	271 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	280 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_Update/ca
      -- CP-element group 277: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_Update/$exit
      -- CP-element group 277: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2437_update_completed_
      -- 
    ca_5825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2437_inst_ack_1, ack => convolution3D_CP_3583_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	271 
    -- CP-element group 278: successors 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_Sample/ra
      -- CP-element group 278: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_Sample/$exit
      -- CP-element group 278: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_sample_completed_
      -- 
    ra_5834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2441_inst_ack_0, ack => convolution3D_CP_3583_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	271 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_Update/$exit
      -- CP-element group 279: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_Update/ca
      -- CP-element group 279: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/type_cast_2441_update_completed_
      -- 
    ca_5839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2441_inst_ack_1, ack => convolution3D_CP_3583_elements(279)); -- 
    -- CP-element group 280:  join  transition  output  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: 	277 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_Sample/crr
      -- CP-element group 280: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_sample_start_
      -- 
    crr_5847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(280), ack => call_stmt_2454_call_req_0); -- 
    convolution3D_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(279) & convolution3D_CP_3583_elements(277);
      gj_convolution3D_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_Sample/cra
      -- CP-element group 281: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_sample_completed_
      -- 
    cra_5848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2454_call_ack_0, ack => convolution3D_CP_3583_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	271 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_Update/cca
      -- CP-element group 282: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/call_stmt_2454_update_completed_
      -- 
    cca_5853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2454_call_ack_1, ack => convolution3D_CP_3583_elements(282)); -- 
    -- CP-element group 283:  join  fork  transition  place  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: 	275 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	297 
    -- CP-element group 283: 	298 
    -- CP-element group 283: 	299 
    -- CP-element group 283: 	284 
    -- CP-element group 283: 	285 
    -- CP-element group 283: 	286 
    -- CP-element group 283: 	287 
    -- CP-element group 283: 	291 
    -- CP-element group 283: 	292 
    -- CP-element group 283: 	293 
    -- CP-element group 283: 	288 
    -- CP-element group 283: 	289 
    -- CP-element group 283: 	290 
    -- CP-element group 283: 	294 
    -- CP-element group 283: 	295 
    -- CP-element group 283: 	296 
    -- CP-element group 283:  members (52) 
      -- CP-element group 283: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454__exit__
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553__entry__
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_1215/call_stmt_2424_to_call_stmt_2454/$exit
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_update_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_update_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_update_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_update_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_update_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_update_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_update_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_update_start_
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_Update/cr
      -- 
    rr_5864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2458_inst_req_0); -- 
    rr_5878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2468_inst_req_0); -- 
    cr_5883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2468_inst_req_1); -- 
    cr_5869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2458_inst_req_1); -- 
    rr_5892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2478_inst_req_0); -- 
    cr_5897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2478_inst_req_1); -- 
    rr_5906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2488_inst_req_0); -- 
    cr_5911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2488_inst_req_1); -- 
    rr_5920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2498_inst_req_0); -- 
    cr_5925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2498_inst_req_1); -- 
    rr_5934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2508_inst_req_0); -- 
    cr_5939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2508_inst_req_1); -- 
    rr_5948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2518_inst_req_0); -- 
    cr_5953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2518_inst_req_1); -- 
    rr_5962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2528_inst_req_0); -- 
    cr_5967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(283), ack => type_cast_2528_inst_req_1); -- 
    convolution3D_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(282) & convolution3D_CP_3583_elements(275);
      gj_convolution3D_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_Sample/ra
      -- 
    ra_5865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2458_inst_ack_0, ack => convolution3D_CP_3583_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	283 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	320 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_Update/ca
      -- CP-element group 285: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2458_Update/$exit
      -- 
    ca_5870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2458_inst_ack_1, ack => convolution3D_CP_3583_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	283 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_sample_completed_
      -- CP-element group 286: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_Sample/ra
      -- CP-element group 286: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_Sample/$exit
      -- 
    ra_5879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2468_inst_ack_0, ack => convolution3D_CP_3583_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	283 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	317 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_update_completed_
      -- CP-element group 287: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2468_Update/$exit
      -- 
    ca_5884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2468_inst_ack_1, ack => convolution3D_CP_3583_elements(287)); -- 
    -- CP-element group 288:  transition  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	283 
    -- CP-element group 288: successors 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_Sample/ra
      -- 
    ra_5893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2478_inst_ack_0, ack => convolution3D_CP_3583_elements(288)); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	283 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	314 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2478_Update/ca
      -- 
    ca_5898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2478_inst_ack_1, ack => convolution3D_CP_3583_elements(289)); -- 
    -- CP-element group 290:  transition  input  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	283 
    -- CP-element group 290: successors 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_sample_completed_
      -- CP-element group 290: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_Sample/$exit
      -- CP-element group 290: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_Sample/ra
      -- 
    ra_5907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2488_inst_ack_0, ack => convolution3D_CP_3583_elements(290)); -- 
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	283 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	311 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_update_completed_
      -- CP-element group 291: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_Update/$exit
      -- CP-element group 291: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2488_Update/ca
      -- 
    ca_5912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2488_inst_ack_1, ack => convolution3D_CP_3583_elements(291)); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	283 
    -- CP-element group 292: successors 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_sample_completed_
      -- CP-element group 292: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_Sample/ra
      -- 
    ra_5921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2498_inst_ack_0, ack => convolution3D_CP_3583_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	283 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	308 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2498_Update/ca
      -- 
    ca_5926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2498_inst_ack_1, ack => convolution3D_CP_3583_elements(293)); -- 
    -- CP-element group 294:  transition  input  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	283 
    -- CP-element group 294: successors 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_sample_completed_
      -- CP-element group 294: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_Sample/$exit
      -- CP-element group 294: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_Sample/ra
      -- 
    ra_5935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_0, ack => convolution3D_CP_3583_elements(294)); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	283 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	305 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_update_completed_
      -- CP-element group 295: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2508_Update/ca
      -- 
    ca_5940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2508_inst_ack_1, ack => convolution3D_CP_3583_elements(295)); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	283 
    -- CP-element group 296: successors 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_sample_completed_
      -- CP-element group 296: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_Sample/ra
      -- 
    ra_5949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2518_inst_ack_0, ack => convolution3D_CP_3583_elements(296)); -- 
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	283 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	302 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_update_completed_
      -- CP-element group 297: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2518_Update/ca
      -- 
    ca_5954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2518_inst_ack_1, ack => convolution3D_CP_3583_elements(297)); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	283 
    -- CP-element group 298: successors 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_sample_completed_
      -- CP-element group 298: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_Sample/$exit
      -- CP-element group 298: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_Sample/ra
      -- 
    ra_5963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2528_inst_ack_0, ack => convolution3D_CP_3583_elements(298)); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	283 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_update_completed_
      -- CP-element group 299: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_Update/$exit
      -- CP-element group 299: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/type_cast_2528_Update/ca
      -- CP-element group 299: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_sample_start_
      -- CP-element group 299: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_Sample/$entry
      -- CP-element group 299: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_Sample/req
      -- 
    ca_5968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2528_inst_ack_1, ack => convolution3D_CP_3583_elements(299)); -- 
    req_5976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(299), ack => WPIPE_maxpool_output_pipe_2530_inst_req_0); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_update_start_
      -- CP-element group 300: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_Sample/ack
      -- CP-element group 300: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_Update/req
      -- 
    ack_5977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2530_inst_ack_0, ack => convolution3D_CP_3583_elements(300)); -- 
    req_5981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(300), ack => WPIPE_maxpool_output_pipe_2530_inst_req_1); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2530_Update/ack
      -- 
    ack_5982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2530_inst_ack_1, ack => convolution3D_CP_3583_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	297 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_Sample/req
      -- 
    req_5990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(302), ack => WPIPE_maxpool_output_pipe_2533_inst_req_0); -- 
    convolution3D_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(297) & convolution3D_CP_3583_elements(301);
      gj_convolution3D_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_update_start_
      -- CP-element group 303: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_Update/req
      -- 
    ack_5991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2533_inst_ack_0, ack => convolution3D_CP_3583_elements(303)); -- 
    req_5995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(303), ack => WPIPE_maxpool_output_pipe_2533_inst_req_1); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2533_Update/ack
      -- 
    ack_5996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2533_inst_ack_1, ack => convolution3D_CP_3583_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	295 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_Sample/req
      -- 
    req_6004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(305), ack => WPIPE_maxpool_output_pipe_2536_inst_req_0); -- 
    convolution3D_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(295) & convolution3D_CP_3583_elements(304);
      gj_convolution3D_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_sample_completed_
      -- CP-element group 306: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_update_start_
      -- CP-element group 306: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_Sample/ack
      -- CP-element group 306: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_Update/req
      -- 
    ack_6005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2536_inst_ack_0, ack => convolution3D_CP_3583_elements(306)); -- 
    req_6009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(306), ack => WPIPE_maxpool_output_pipe_2536_inst_req_1); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_update_completed_
      -- CP-element group 307: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2536_Update/ack
      -- 
    ack_6010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2536_inst_ack_1, ack => convolution3D_CP_3583_elements(307)); -- 
    -- CP-element group 308:  join  transition  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	293 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_Sample/req
      -- 
    req_6018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(308), ack => WPIPE_maxpool_output_pipe_2539_inst_req_0); -- 
    convolution3D_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(293) & convolution3D_CP_3583_elements(307);
      gj_convolution3D_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_update_start_
      -- CP-element group 309: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_Update/req
      -- 
    ack_6019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2539_inst_ack_0, ack => convolution3D_CP_3583_elements(309)); -- 
    req_6023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(309), ack => WPIPE_maxpool_output_pipe_2539_inst_req_1); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2539_Update/ack
      -- 
    ack_6024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2539_inst_ack_1, ack => convolution3D_CP_3583_elements(310)); -- 
    -- CP-element group 311:  join  transition  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	291 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_sample_start_
      -- CP-element group 311: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_Sample/req
      -- 
    req_6032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(311), ack => WPIPE_maxpool_output_pipe_2542_inst_req_0); -- 
    convolution3D_cp_element_group_311: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_311"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(291) & convolution3D_CP_3583_elements(310);
      gj_convolution3D_cp_element_group_311 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(311), clk => clk, reset => reset); --
    end block;
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_sample_completed_
      -- CP-element group 312: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_update_start_
      -- CP-element group 312: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_Sample/ack
      -- CP-element group 312: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_Update/req
      -- 
    ack_6033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2542_inst_ack_0, ack => convolution3D_CP_3583_elements(312)); -- 
    req_6037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(312), ack => WPIPE_maxpool_output_pipe_2542_inst_req_1); -- 
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_update_completed_
      -- CP-element group 313: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2542_Update/ack
      -- 
    ack_6038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2542_inst_ack_1, ack => convolution3D_CP_3583_elements(313)); -- 
    -- CP-element group 314:  join  transition  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	289 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_sample_start_
      -- CP-element group 314: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_Sample/$entry
      -- CP-element group 314: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_Sample/req
      -- 
    req_6046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(314), ack => WPIPE_maxpool_output_pipe_2545_inst_req_0); -- 
    convolution3D_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(289) & convolution3D_CP_3583_elements(313);
      gj_convolution3D_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  transition  input  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (6) 
      -- CP-element group 315: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_update_start_
      -- CP-element group 315: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_Sample/ack
      -- CP-element group 315: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_Update/req
      -- 
    ack_6047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2545_inst_ack_0, ack => convolution3D_CP_3583_elements(315)); -- 
    req_6051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(315), ack => WPIPE_maxpool_output_pipe_2545_inst_req_1); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2545_Update/ack
      -- 
    ack_6052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2545_inst_ack_1, ack => convolution3D_CP_3583_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	287 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_Sample/req
      -- 
    req_6060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(317), ack => WPIPE_maxpool_output_pipe_2548_inst_req_0); -- 
    convolution3D_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(287) & convolution3D_CP_3583_elements(316);
      gj_convolution3D_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_update_start_
      -- CP-element group 318: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_Update/req
      -- 
    ack_6061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2548_inst_ack_0, ack => convolution3D_CP_3583_elements(318)); -- 
    req_6065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(318), ack => WPIPE_maxpool_output_pipe_2548_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2548_Update/ack
      -- 
    ack_6066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2548_inst_ack_1, ack => convolution3D_CP_3583_elements(319)); -- 
    -- CP-element group 320:  join  transition  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	285 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_sample_start_
      -- CP-element group 320: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_Sample/$entry
      -- CP-element group 320: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_Sample/req
      -- 
    req_6074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(320), ack => WPIPE_maxpool_output_pipe_2551_inst_req_0); -- 
    convolution3D_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(285) & convolution3D_CP_3583_elements(319);
      gj_convolution3D_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  transition  input  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (6) 
      -- CP-element group 321: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_sample_completed_
      -- CP-element group 321: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_update_start_
      -- CP-element group 321: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_Sample/ack
      -- CP-element group 321: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_Update/$entry
      -- CP-element group 321: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_Update/req
      -- 
    ack_6075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2551_inst_ack_0, ack => convolution3D_CP_3583_elements(321)); -- 
    req_6079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(321), ack => WPIPE_maxpool_output_pipe_2551_inst_req_1); -- 
    -- CP-element group 322:  transition  place  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322:  members (16) 
      -- CP-element group 322: 	 branch_block_stmt_1215/return__
      -- CP-element group 322: 	 branch_block_stmt_1215/merge_stmt_2555__exit__
      -- CP-element group 322: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553__exit__
      -- CP-element group 322: 	 branch_block_stmt_1215/$exit
      -- CP-element group 322: 	 branch_block_stmt_1215/branch_block_stmt_1215__exit__
      -- CP-element group 322: 	 $exit
      -- CP-element group 322: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/$exit
      -- CP-element group 322: 	 branch_block_stmt_1215/merge_stmt_2555_PhiAck/dummy
      -- CP-element group 322: 	 branch_block_stmt_1215/merge_stmt_2555_PhiAck/$exit
      -- CP-element group 322: 	 branch_block_stmt_1215/merge_stmt_2555_PhiAck/$entry
      -- CP-element group 322: 	 branch_block_stmt_1215/return___PhiReq/$exit
      -- CP-element group 322: 	 branch_block_stmt_1215/return___PhiReq/$entry
      -- CP-element group 322: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_update_completed_
      -- CP-element group 322: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_1215/assign_stmt_2459_to_assign_stmt_2553/WPIPE_maxpool_output_pipe_2551_Update/ack
      -- CP-element group 322: 	 branch_block_stmt_1215/merge_stmt_2555_PhiReqMerge
      -- 
    ack_6080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2551_inst_ack_1, ack => convolution3D_CP_3583_elements(322)); -- 
    -- CP-element group 323:  transition  output  delay-element  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	80 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	327 
    -- CP-element group 323:  members (5) 
      -- CP-element group 323: 	 branch_block_stmt_1215/bbx_xnph370_forx_xbody_PhiReq/$exit
      -- CP-element group 323: 	 branch_block_stmt_1215/bbx_xnph370_forx_xbody_PhiReq/phi_stmt_1524/$exit
      -- CP-element group 323: 	 branch_block_stmt_1215/bbx_xnph370_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/$exit
      -- CP-element group 323: 	 branch_block_stmt_1215/bbx_xnph370_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1528_konst_delay_trans
      -- CP-element group 323: 	 branch_block_stmt_1215/bbx_xnph370_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_req
      -- 
    phi_stmt_1524_req_6103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1524_req_6103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(323), ack => phi_stmt_1524_req_0); -- 
    -- Element group convolution3D_CP_3583_elements(323) is a control-delay.
    cp_element_323_delay: control_delay_element  generic map(name => " 323_delay", delay_value => 1)  port map(req => convolution3D_CP_3583_elements(80), ack => convolution3D_CP_3583_elements(323), clk => clk, reset =>reset);
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	122 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (2) 
      -- CP-element group 324: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/SplitProtocol/Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/SplitProtocol/Sample/ra
      -- 
    ra_6123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1530_inst_ack_0, ack => convolution3D_CP_3583_elements(324)); -- 
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	122 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (2) 
      -- CP-element group 325: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/SplitProtocol/Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/SplitProtocol/Update/ca
      -- 
    ca_6128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1530_inst_ack_1, ack => convolution3D_CP_3583_elements(325)); -- 
    -- CP-element group 326:  join  transition  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 326: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/$exit
      -- CP-element group 326: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/$exit
      -- CP-element group 326: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/$exit
      -- CP-element group 326: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_sources/type_cast_1530/SplitProtocol/$exit
      -- CP-element group 326: 	 branch_block_stmt_1215/forx_xbody_forx_xbody_PhiReq/phi_stmt_1524/phi_stmt_1524_req
      -- 
    phi_stmt_1524_req_6129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1524_req_6129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(326), ack => phi_stmt_1524_req_1); -- 
    convolution3D_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(324) & convolution3D_CP_3583_elements(325);
      gj_convolution3D_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  merge  transition  place  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	323 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (2) 
      -- CP-element group 327: 	 branch_block_stmt_1215/merge_stmt_1523_PhiReqMerge
      -- CP-element group 327: 	 branch_block_stmt_1215/merge_stmt_1523_PhiAck/$entry
      -- 
    convolution3D_CP_3583_elements(327) <= OrReduce(convolution3D_CP_3583_elements(323) & convolution3D_CP_3583_elements(326));
    -- CP-element group 328:  fork  transition  place  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	96 
    -- CP-element group 328: 	104 
    -- CP-element group 328: 	112 
    -- CP-element group 328: 	108 
    -- CP-element group 328: 	100 
    -- CP-element group 328: 	116 
    -- CP-element group 328: 	119 
    -- CP-element group 328: 	81 
    -- CP-element group 328: 	82 
    -- CP-element group 328: 	84 
    -- CP-element group 328: 	85 
    -- CP-element group 328: 	88 
    -- CP-element group 328: 	92 
    -- CP-element group 328:  members (56) 
      -- CP-element group 328: 	 branch_block_stmt_1215/merge_stmt_1523__exit__
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686__entry__
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_update_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_resized_1
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_scaled_1
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_computed_1
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_resize_1/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_resize_1/$exit
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_resize_1/index_resize_req
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_resize_1/index_resize_ack
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_scale_1/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_scale_1/$exit
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_scale_1/scale_rename_req
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_index_scale_1/scale_rename_ack
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_final_index_sum_regn_update_start
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_final_index_sum_regn_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_final_index_sum_regn_Sample/req
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_final_index_sum_regn_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/array_obj_ref_1536_final_index_sum_regn_Update/req
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_complete/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/addr_of_1537_complete/req
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/RPIPE_maxpool_input_pipe_1540_Sample/rr
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_update_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1544_Update/cr
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_update_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1557_Update/cr
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_update_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1575_Update/cr
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_update_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1593_Update/cr
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_update_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1611_Update/cr
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_update_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1629_Update/cr
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_update_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1647_Update/cr
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_update_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/type_cast_1665_Update/cr
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_update_start_
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Update/word_access_complete/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Update/word_access_complete/word_0/$entry
      -- CP-element group 328: 	 branch_block_stmt_1215/assign_stmt_1538_to_assign_stmt_1686/ptr_deref_1673_Update/word_access_complete/word_0/cr
      -- CP-element group 328: 	 branch_block_stmt_1215/merge_stmt_1523_PhiAck/$exit
      -- CP-element group 328: 	 branch_block_stmt_1215/merge_stmt_1523_PhiAck/phi_stmt_1524_ack
      -- 
    phi_stmt_1524_ack_6134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1524_ack_0, ack => convolution3D_CP_3583_elements(328)); -- 
    req_4263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => array_obj_ref_1536_index_offset_req_0); -- 
    req_4268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => array_obj_ref_1536_index_offset_req_1); -- 
    req_4283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => addr_of_1537_final_reg_req_1); -- 
    rr_4292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => RPIPE_maxpool_input_pipe_1540_inst_req_0); -- 
    cr_4311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => type_cast_1544_inst_req_1); -- 
    cr_4339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => type_cast_1557_inst_req_1); -- 
    cr_4367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => type_cast_1575_inst_req_1); -- 
    cr_4395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => type_cast_1593_inst_req_1); -- 
    cr_4423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => type_cast_1611_inst_req_1); -- 
    cr_4451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => type_cast_1629_inst_req_1); -- 
    cr_4479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => type_cast_1647_inst_req_1); -- 
    cr_4507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => type_cast_1665_inst_req_1); -- 
    cr_4557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(328), ack => ptr_deref_1673_store_0_req_1); -- 
    -- CP-element group 329:  transition  output  delay-element  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	73 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	333 
    -- CP-element group 329:  members (5) 
      -- CP-element group 329: 	 branch_block_stmt_1215/entry_forx_xend_PhiReq/$exit
      -- CP-element group 329: 	 branch_block_stmt_1215/entry_forx_xend_PhiReq/phi_stmt_1707/$exit
      -- CP-element group 329: 	 branch_block_stmt_1215/entry_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/$exit
      -- CP-element group 329: 	 branch_block_stmt_1215/entry_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1713_konst_delay_trans
      -- CP-element group 329: 	 branch_block_stmt_1215/entry_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_req
      -- 
    phi_stmt_1707_req_6157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1707_req_6157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(329), ack => phi_stmt_1707_req_1); -- 
    -- Element group convolution3D_CP_3583_elements(329) is a control-delay.
    cp_element_329_delay: control_delay_element  generic map(name => " 329_delay", delay_value => 1)  port map(req => convolution3D_CP_3583_elements(73), ack => convolution3D_CP_3583_elements(329), clk => clk, reset =>reset);
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	124 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	332 
    -- CP-element group 330:  members (2) 
      -- CP-element group 330: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Sample/$exit
      -- CP-element group 330: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Sample/ra
      -- 
    ra_6177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1710_inst_ack_0, ack => convolution3D_CP_3583_elements(330)); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	124 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (2) 
      -- CP-element group 331: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Update/$exit
      -- CP-element group 331: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/Update/ca
      -- 
    ca_6182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1710_inst_ack_1, ack => convolution3D_CP_3583_elements(331)); -- 
    -- CP-element group 332:  join  transition  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: 	330 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 332: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/$exit
      -- CP-element group 332: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/$exit
      -- CP-element group 332: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/$exit
      -- CP-element group 332: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_sources/type_cast_1710/SplitProtocol/$exit
      -- CP-element group 332: 	 branch_block_stmt_1215/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1707/phi_stmt_1707_req
      -- 
    phi_stmt_1707_req_6183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1707_req_6183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(332), ack => phi_stmt_1707_req_0); -- 
    convolution3D_cp_element_group_332: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_332"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(331) & convolution3D_CP_3583_elements(330);
      gj_convolution3D_cp_element_group_332 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(332), clk => clk, reset => reset); --
    end block;
    -- CP-element group 333:  merge  transition  place  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: 	329 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (2) 
      -- CP-element group 333: 	 branch_block_stmt_1215/merge_stmt_1706_PhiReqMerge
      -- CP-element group 333: 	 branch_block_stmt_1215/merge_stmt_1706_PhiAck/$entry
      -- 
    convolution3D_CP_3583_elements(333) <= OrReduce(convolution3D_CP_3583_elements(332) & convolution3D_CP_3583_elements(329));
    -- CP-element group 334:  branch  transition  place  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	125 
    -- CP-element group 334: 	126 
    -- CP-element group 334:  members (15) 
      -- CP-element group 334: 	 branch_block_stmt_1215/assign_stmt_1720_to_assign_stmt_1726__entry__
      -- CP-element group 334: 	 branch_block_stmt_1215/merge_stmt_1706__exit__
      -- CP-element group 334: 	 branch_block_stmt_1215/assign_stmt_1720_to_assign_stmt_1726__exit__
      -- CP-element group 334: 	 branch_block_stmt_1215/R_tobool_1728_place
      -- CP-element group 334: 	 branch_block_stmt_1215/if_stmt_1727_else_link/$entry
      -- CP-element group 334: 	 branch_block_stmt_1215/if_stmt_1727__entry__
      -- CP-element group 334: 	 branch_block_stmt_1215/if_stmt_1727_if_link/$entry
      -- CP-element group 334: 	 branch_block_stmt_1215/assign_stmt_1720_to_assign_stmt_1726/$entry
      -- CP-element group 334: 	 branch_block_stmt_1215/assign_stmt_1720_to_assign_stmt_1726/$exit
      -- CP-element group 334: 	 branch_block_stmt_1215/if_stmt_1727_dead_link/$entry
      -- CP-element group 334: 	 branch_block_stmt_1215/if_stmt_1727_eval_test/$entry
      -- CP-element group 334: 	 branch_block_stmt_1215/if_stmt_1727_eval_test/$exit
      -- CP-element group 334: 	 branch_block_stmt_1215/if_stmt_1727_eval_test/branch_req
      -- CP-element group 334: 	 branch_block_stmt_1215/merge_stmt_1706_PhiAck/$exit
      -- CP-element group 334: 	 branch_block_stmt_1215/merge_stmt_1706_PhiAck/phi_stmt_1707_ack
      -- 
    phi_stmt_1707_ack_6188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1707_ack_0, ack => convolution3D_CP_3583_elements(334)); -- 
    branch_req_4605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(334), ack => if_stmt_1727_branch_req_0); -- 
    -- CP-element group 335:  transition  input  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	141 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (2) 
      -- CP-element group 335: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Sample/ra
      -- 
    ra_6220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1773_inst_ack_0, ack => convolution3D_CP_3583_elements(335)); -- 
    -- CP-element group 336:  transition  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	141 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (2) 
      -- CP-element group 336: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/Update/ca
      -- 
    ca_6225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1773_inst_ack_1, ack => convolution3D_CP_3583_elements(336)); -- 
    -- CP-element group 337:  join  transition  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	341 
    -- CP-element group 337:  members (5) 
      -- CP-element group 337: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/$exit
      -- CP-element group 337: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/$exit
      -- CP-element group 337: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/$exit
      -- CP-element group 337: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1773/SplitProtocol/$exit
      -- CP-element group 337: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_req
      -- 
    phi_stmt_1770_req_6226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1770_req_6226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(337), ack => phi_stmt_1770_req_0); -- 
    convolution3D_cp_element_group_337: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_337"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(335) & convolution3D_CP_3583_elements(336);
      gj_convolution3D_cp_element_group_337 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(337), clk => clk, reset => reset); --
    end block;
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	141 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (2) 
      -- CP-element group 338: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/SplitProtocol/Sample/$exit
      -- CP-element group 338: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/SplitProtocol/Sample/ra
      -- 
    ra_6243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1766_inst_ack_0, ack => convolution3D_CP_3583_elements(338)); -- 
    -- CP-element group 339:  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	141 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (2) 
      -- CP-element group 339: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/SplitProtocol/Update/$exit
      -- CP-element group 339: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/SplitProtocol/Update/ca
      -- 
    ca_6248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1766_inst_ack_1, ack => convolution3D_CP_3583_elements(339)); -- 
    -- CP-element group 340:  join  transition  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (5) 
      -- CP-element group 340: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/$exit
      -- CP-element group 340: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/$exit
      -- CP-element group 340: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/$exit
      -- CP-element group 340: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1766/SplitProtocol/$exit
      -- CP-element group 340: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_req
      -- 
    phi_stmt_1763_req_6249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1763_req_6249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(340), ack => phi_stmt_1763_req_0); -- 
    convolution3D_cp_element_group_340: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_340"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(338) & convolution3D_CP_3583_elements(339);
      gj_convolution3D_cp_element_group_340 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(340), clk => clk, reset => reset); --
    end block;
    -- CP-element group 341:  join  transition  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	337 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	345 
    -- CP-element group 341:  members (1) 
      -- CP-element group 341: 	 branch_block_stmt_1215/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_341: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_341"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(337) & convolution3D_CP_3583_elements(340);
      gj_convolution3D_cp_element_group_341 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(341), clk => clk, reset => reset); --
    end block;
    -- CP-element group 342:  transition  output  delay-element  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	135 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (4) 
      -- CP-element group 342: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1770/$exit
      -- CP-element group 342: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/$exit
      -- CP-element group 342: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_sources/type_cast_1776_konst_delay_trans
      -- CP-element group 342: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1770/phi_stmt_1770_req
      -- 
    phi_stmt_1770_req_6260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1770_req_6260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(342), ack => phi_stmt_1770_req_1); -- 
    -- Element group convolution3D_CP_3583_elements(342) is a control-delay.
    cp_element_342_delay: control_delay_element  generic map(name => " 342_delay", delay_value => 1)  port map(req => convolution3D_CP_3583_elements(135), ack => convolution3D_CP_3583_elements(342), clk => clk, reset =>reset);
    -- CP-element group 343:  transition  output  delay-element  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	135 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (4) 
      -- CP-element group 343: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1763/$exit
      -- CP-element group 343: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/$exit
      -- CP-element group 343: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_sources/type_cast_1769_konst_delay_trans
      -- CP-element group 343: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1763/phi_stmt_1763_req
      -- 
    phi_stmt_1763_req_6268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1763_req_6268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(343), ack => phi_stmt_1763_req_1); -- 
    -- Element group convolution3D_CP_3583_elements(343) is a control-delay.
    cp_element_343_delay: control_delay_element  generic map(name => " 343_delay", delay_value => 1)  port map(req => convolution3D_CP_3583_elements(135), ack => convolution3D_CP_3583_elements(343), clk => clk, reset =>reset);
    -- CP-element group 344:  join  transition  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (1) 
      -- CP-element group 344: 	 branch_block_stmt_1215/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_344: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_344"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(342) & convolution3D_CP_3583_elements(343);
      gj_convolution3D_cp_element_group_344 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(344), clk => clk, reset => reset); --
    end block;
    -- CP-element group 345:  merge  fork  transition  place  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	341 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (2) 
      -- CP-element group 345: 	 branch_block_stmt_1215/merge_stmt_1762_PhiReqMerge
      -- CP-element group 345: 	 branch_block_stmt_1215/merge_stmt_1762_PhiAck/$entry
      -- 
    convolution3D_CP_3583_elements(345) <= OrReduce(convolution3D_CP_3583_elements(341) & convolution3D_CP_3583_elements(344));
    -- CP-element group 346:  transition  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (1) 
      -- CP-element group 346: 	 branch_block_stmt_1215/merge_stmt_1762_PhiAck/phi_stmt_1763_ack
      -- 
    phi_stmt_1763_ack_6273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1763_ack_0, ack => convolution3D_CP_3583_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (1) 
      -- CP-element group 347: 	 branch_block_stmt_1215/merge_stmt_1762_PhiAck/phi_stmt_1770_ack
      -- 
    phi_stmt_1770_ack_6274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1770_ack_0, ack => convolution3D_CP_3583_elements(347)); -- 
    -- CP-element group 348:  join  fork  transition  place  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	136 
    -- CP-element group 348: 	139 
    -- CP-element group 348:  members (10) 
      -- CP-element group 348: 	 branch_block_stmt_1215/merge_stmt_1762__exit__
      -- CP-element group 348: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806__entry__
      -- CP-element group 348: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_Update/cr
      -- CP-element group 348: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/type_cast_1783_update_start_
      -- CP-element group 348: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_Sample/rr
      -- CP-element group 348: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_Sample/$entry
      -- CP-element group 348: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/RPIPE_maxpool_input_pipe_1779_sample_start_
      -- CP-element group 348: 	 branch_block_stmt_1215/assign_stmt_1780_to_assign_stmt_1806/$entry
      -- CP-element group 348: 	 branch_block_stmt_1215/merge_stmt_1762_PhiAck/$exit
      -- 
    cr_4705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(348), ack => type_cast_1783_inst_req_1); -- 
    rr_4686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(348), ack => RPIPE_maxpool_input_pipe_1779_inst_req_0); -- 
    convolution3D_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(346) & convolution3D_CP_3583_elements(347);
      gj_convolution3D_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	140 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	351 
    -- CP-element group 349:  members (2) 
      -- CP-element group 349: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/SplitProtocol/Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/SplitProtocol/Sample/ra
      -- 
    ra_6298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1817_inst_ack_0, ack => convolution3D_CP_3583_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	140 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (2) 
      -- CP-element group 350: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/SplitProtocol/Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/SplitProtocol/Update/ca
      -- 
    ca_6303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1817_inst_ack_1, ack => convolution3D_CP_3583_elements(350)); -- 
    -- CP-element group 351:  join  transition  place  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	349 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (8) 
      -- CP-element group 351: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 351: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/$exit
      -- CP-element group 351: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/$exit
      -- CP-element group 351: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/$exit
      -- CP-element group 351: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_sources/type_cast_1817/SplitProtocol/$exit
      -- CP-element group 351: 	 branch_block_stmt_1215/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1814/phi_stmt_1814_req
      -- CP-element group 351: 	 branch_block_stmt_1215/merge_stmt_1813_PhiReqMerge
      -- CP-element group 351: 	 branch_block_stmt_1215/merge_stmt_1813_PhiAck/$entry
      -- 
    phi_stmt_1814_req_6304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1814_req_6304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(351), ack => phi_stmt_1814_req_0); -- 
    convolution3D_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(349) & convolution3D_CP_3583_elements(350);
      gj_convolution3D_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	150 
    -- CP-element group 352: 	144 
    -- CP-element group 352: 	145 
    -- CP-element group 352: 	147 
    -- CP-element group 352: 	142 
    -- CP-element group 352: 	143 
    -- CP-element group 352:  members (35) 
      -- CP-element group 352: 	 branch_block_stmt_1215/merge_stmt_1813__exit__
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856__entry__
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_Update/cr
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_update_start_
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Update/word_access_complete/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_Sample/rr
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_update_start_
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_update_start_
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/type_cast_1821_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_complete/req
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/addr_of_1851_complete/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_final_index_sum_regn_Update/req
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_final_index_sum_regn_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_final_index_sum_regn_Sample/req
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_final_index_sum_regn_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_final_index_sum_regn_update_start
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_scale_1/scale_rename_ack
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Update/word_access_complete/word_0/cr
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/ptr_deref_1854_Update/word_access_complete/word_0/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_scale_1/scale_rename_req
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_scale_1/$exit
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_scale_1/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_resize_1/index_resize_ack
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_resize_1/index_resize_req
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_resize_1/$exit
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_resize_1/$entry
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_computed_1
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_scaled_1
      -- CP-element group 352: 	 branch_block_stmt_1215/assign_stmt_1822_to_assign_stmt_1856/array_obj_ref_1850_index_resized_1
      -- CP-element group 352: 	 branch_block_stmt_1215/merge_stmt_1813_PhiAck/$exit
      -- CP-element group 352: 	 branch_block_stmt_1215/merge_stmt_1813_PhiAck/phi_stmt_1814_ack
      -- 
    phi_stmt_1814_ack_6309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1814_ack_0, ack => convolution3D_CP_3583_elements(352)); -- 
    cr_4741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(352), ack => type_cast_1821_inst_req_1); -- 
    rr_4736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(352), ack => type_cast_1821_inst_req_0); -- 
    req_4787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(352), ack => addr_of_1851_final_reg_req_1); -- 
    req_4772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(352), ack => array_obj_ref_1850_index_offset_req_1); -- 
    req_4767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(352), ack => array_obj_ref_1850_index_offset_req_0); -- 
    cr_4837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(352), ack => ptr_deref_1854_store_0_req_1); -- 
    -- CP-element group 353:  merge  fork  transition  place  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	151 
    -- CP-element group 353: 	125 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	154 
    -- CP-element group 353: 	155 
    -- CP-element group 353: 	152 
    -- CP-element group 353: 	153 
    -- CP-element group 353: 	156 
    -- CP-element group 353: 	157 
    -- CP-element group 353:  members (25) 
      -- CP-element group 353: 	 branch_block_stmt_1215/merge_stmt_1858__exit__
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_Update/cr
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891__entry__
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_Sample/rr
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_Update/cr
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_update_start_
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_Sample/rr
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1869_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_Update/cr
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_update_start_
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1861_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/$entry
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_Sample/rr
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_update_start_
      -- CP-element group 353: 	 branch_block_stmt_1215/assign_stmt_1862_to_assign_stmt_1891/type_cast_1865_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_1215/merge_stmt_1858_PhiReqMerge
      -- CP-element group 353: 	 branch_block_stmt_1215/merge_stmt_1858_PhiAck/$entry
      -- CP-element group 353: 	 branch_block_stmt_1215/merge_stmt_1858_PhiAck/$exit
      -- CP-element group 353: 	 branch_block_stmt_1215/merge_stmt_1858_PhiAck/dummy
      -- 
    cr_4882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(353), ack => type_cast_1869_inst_req_1); -- 
    rr_4877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(353), ack => type_cast_1869_inst_req_0); -- 
    cr_4854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(353), ack => type_cast_1861_inst_req_1); -- 
    rr_4849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(353), ack => type_cast_1861_inst_req_0); -- 
    cr_4868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(353), ack => type_cast_1865_inst_req_1); -- 
    rr_4863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(353), ack => type_cast_1865_inst_req_0); -- 
    convolution3D_CP_3583_elements(353) <= OrReduce(convolution3D_CP_3583_elements(151) & convolution3D_CP_3583_elements(125));
    -- CP-element group 354:  transition  output  delay-element  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	171 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	358 
    -- CP-element group 354:  members (5) 
      -- CP-element group 354: 	 branch_block_stmt_1215/bbx_xnph_forx_xbody159_PhiReq/$exit
      -- CP-element group 354: 	 branch_block_stmt_1215/bbx_xnph_forx_xbody159_PhiReq/phi_stmt_1979/$exit
      -- CP-element group 354: 	 branch_block_stmt_1215/bbx_xnph_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/$exit
      -- CP-element group 354: 	 branch_block_stmt_1215/bbx_xnph_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1983_konst_delay_trans
      -- CP-element group 354: 	 branch_block_stmt_1215/bbx_xnph_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_req
      -- 
    phi_stmt_1979_req_6343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1979_req_6343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(354), ack => phi_stmt_1979_req_0); -- 
    -- Element group convolution3D_CP_3583_elements(354) is a control-delay.
    cp_element_354_delay: control_delay_element  generic map(name => " 354_delay", delay_value => 1)  port map(req => convolution3D_CP_3583_elements(171), ack => convolution3D_CP_3583_elements(354), clk => clk, reset =>reset);
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	213 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	357 
    -- CP-element group 355:  members (2) 
      -- CP-element group 355: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/SplitProtocol/Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/SplitProtocol/Sample/ra
      -- 
    ra_6363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1985_inst_ack_0, ack => convolution3D_CP_3583_elements(355)); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	213 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (2) 
      -- CP-element group 356: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/SplitProtocol/Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/SplitProtocol/Update/ca
      -- 
    ca_6368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1985_inst_ack_1, ack => convolution3D_CP_3583_elements(356)); -- 
    -- CP-element group 357:  join  transition  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	355 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/$exit
      -- CP-element group 357: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/$exit
      -- CP-element group 357: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/$exit
      -- CP-element group 357: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/$exit
      -- CP-element group 357: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_sources/type_cast_1985/SplitProtocol/$exit
      -- CP-element group 357: 	 branch_block_stmt_1215/forx_xbody159_forx_xbody159_PhiReq/phi_stmt_1979/phi_stmt_1979_req
      -- 
    phi_stmt_1979_req_6369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1979_req_6369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(357), ack => phi_stmt_1979_req_1); -- 
    convolution3D_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(355) & convolution3D_CP_3583_elements(356);
      gj_convolution3D_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  merge  transition  place  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	354 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (2) 
      -- CP-element group 358: 	 branch_block_stmt_1215/merge_stmt_1978_PhiReqMerge
      -- CP-element group 358: 	 branch_block_stmt_1215/merge_stmt_1978_PhiAck/$entry
      -- 
    convolution3D_CP_3583_elements(358) <= OrReduce(convolution3D_CP_3583_elements(354) & convolution3D_CP_3583_elements(357));
    -- CP-element group 359:  fork  transition  place  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	187 
    -- CP-element group 359: 	207 
    -- CP-element group 359: 	176 
    -- CP-element group 359: 	173 
    -- CP-element group 359: 	175 
    -- CP-element group 359: 	199 
    -- CP-element group 359: 	172 
    -- CP-element group 359: 	179 
    -- CP-element group 359: 	210 
    -- CP-element group 359: 	191 
    -- CP-element group 359: 	183 
    -- CP-element group 359: 	195 
    -- CP-element group 359: 	203 
    -- CP-element group 359:  members (56) 
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141__entry__
      -- CP-element group 359: 	 branch_block_stmt_1215/merge_stmt_1978__exit__
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_update_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_resized_1
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_scaled_1
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_computed_1
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_resize_1/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_resize_1/$exit
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_resize_1/index_resize_req
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_resize_1/index_resize_ack
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_scale_1/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_scale_1/$exit
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_scale_1/scale_rename_req
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_index_scale_1/scale_rename_ack
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_final_index_sum_regn_update_start
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_final_index_sum_regn_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_final_index_sum_regn_Sample/req
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_final_index_sum_regn_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/array_obj_ref_1991_final_index_sum_regn_Update/req
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_complete/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/addr_of_1992_complete/req
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_sample_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/RPIPE_maxpool_input_pipe_1995_Sample/rr
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_update_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_1999_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_update_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2012_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_update_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2030_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_update_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2048_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_update_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2066_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_update_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2084_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_update_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2102_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_update_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/type_cast_2120_Update/cr
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_update_start_
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Update/word_access_complete/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Update/word_access_complete/word_0/$entry
      -- CP-element group 359: 	 branch_block_stmt_1215/assign_stmt_1993_to_assign_stmt_2141/ptr_deref_2128_Update/word_access_complete/word_0/cr
      -- CP-element group 359: 	 branch_block_stmt_1215/merge_stmt_1978_PhiAck/$exit
      -- CP-element group 359: 	 branch_block_stmt_1215/merge_stmt_1978_PhiAck/phi_stmt_1979_ack
      -- 
    phi_stmt_1979_ack_6374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1979_ack_0, ack => convolution3D_CP_3583_elements(359)); -- 
    req_5003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => array_obj_ref_1991_index_offset_req_0); -- 
    req_5008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => array_obj_ref_1991_index_offset_req_1); -- 
    req_5023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => addr_of_1992_final_reg_req_1); -- 
    rr_5032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => RPIPE_maxpool_input_pipe_1995_inst_req_0); -- 
    cr_5051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => type_cast_1999_inst_req_1); -- 
    cr_5079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => type_cast_2012_inst_req_1); -- 
    cr_5107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => type_cast_2030_inst_req_1); -- 
    cr_5135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => type_cast_2048_inst_req_1); -- 
    cr_5163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => type_cast_2066_inst_req_1); -- 
    cr_5191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => type_cast_2084_inst_req_1); -- 
    cr_5219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => type_cast_2102_inst_req_1); -- 
    cr_5247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => type_cast_2120_inst_req_1); -- 
    cr_5297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(359), ack => ptr_deref_2128_store_0_req_1); -- 
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	215 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	362 
    -- CP-element group 360:  members (2) 
      -- CP-element group 360: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/SplitProtocol/Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/SplitProtocol/Sample/ra
      -- 
    ra_6406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2165_inst_ack_0, ack => convolution3D_CP_3583_elements(360)); -- 
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	215 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (2) 
      -- CP-element group 361: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/SplitProtocol/Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/SplitProtocol/Update/ca
      -- 
    ca_6411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2165_inst_ack_1, ack => convolution3D_CP_3583_elements(361)); -- 
    -- CP-element group 362:  join  transition  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	360 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/$exit
      -- CP-element group 362: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/$exit
      -- CP-element group 362: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/$exit
      -- CP-element group 362: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/$exit
      -- CP-element group 362: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2165/SplitProtocol/$exit
      -- CP-element group 362: 	 branch_block_stmt_1215/forx_xcond153x_xforx_xend211_crit_edge_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_req
      -- 
    phi_stmt_2162_req_6412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2162_req_6412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(362), ack => phi_stmt_2162_req_0); -- 
    convolution3D_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(360) & convolution3D_CP_3583_elements(361);
      gj_convolution3D_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  transition  output  delay-element  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	160 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (5) 
      -- CP-element group 363: 	 branch_block_stmt_1215/ifx_xend_forx_xend211_PhiReq/$exit
      -- CP-element group 363: 	 branch_block_stmt_1215/ifx_xend_forx_xend211_PhiReq/phi_stmt_2162/$exit
      -- CP-element group 363: 	 branch_block_stmt_1215/ifx_xend_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/$exit
      -- CP-element group 363: 	 branch_block_stmt_1215/ifx_xend_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_sources/type_cast_2168_konst_delay_trans
      -- CP-element group 363: 	 branch_block_stmt_1215/ifx_xend_forx_xend211_PhiReq/phi_stmt_2162/phi_stmt_2162_req
      -- 
    phi_stmt_2162_req_6423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2162_req_6423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(363), ack => phi_stmt_2162_req_1); -- 
    -- Element group convolution3D_CP_3583_elements(363) is a control-delay.
    cp_element_363_delay: control_delay_element  generic map(name => " 363_delay", delay_value => 1)  port map(req => convolution3D_CP_3583_elements(160), ack => convolution3D_CP_3583_elements(363), clk => clk, reset =>reset);
    -- CP-element group 364:  merge  transition  place  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (2) 
      -- CP-element group 364: 	 branch_block_stmt_1215/merge_stmt_2161_PhiReqMerge
      -- CP-element group 364: 	 branch_block_stmt_1215/merge_stmt_2161_PhiAck/$entry
      -- 
    convolution3D_CP_3583_elements(364) <= OrReduce(convolution3D_CP_3583_elements(363) & convolution3D_CP_3583_elements(362));
    -- CP-element group 365:  branch  transition  place  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	216 
    -- CP-element group 365: 	217 
    -- CP-element group 365:  members (15) 
      -- CP-element group 365: 	 branch_block_stmt_1215/assign_stmt_2175_to_assign_stmt_2181__exit__
      -- CP-element group 365: 	 branch_block_stmt_1215/merge_stmt_2161__exit__
      -- CP-element group 365: 	 branch_block_stmt_1215/assign_stmt_2175_to_assign_stmt_2181__entry__
      -- CP-element group 365: 	 branch_block_stmt_1215/if_stmt_2182__entry__
      -- CP-element group 365: 	 branch_block_stmt_1215/assign_stmt_2175_to_assign_stmt_2181/$entry
      -- CP-element group 365: 	 branch_block_stmt_1215/assign_stmt_2175_to_assign_stmt_2181/$exit
      -- CP-element group 365: 	 branch_block_stmt_1215/if_stmt_2182_dead_link/$entry
      -- CP-element group 365: 	 branch_block_stmt_1215/if_stmt_2182_eval_test/$entry
      -- CP-element group 365: 	 branch_block_stmt_1215/if_stmt_2182_eval_test/$exit
      -- CP-element group 365: 	 branch_block_stmt_1215/if_stmt_2182_eval_test/branch_req
      -- CP-element group 365: 	 branch_block_stmt_1215/R_tobool214_2183_place
      -- CP-element group 365: 	 branch_block_stmt_1215/if_stmt_2182_if_link/$entry
      -- CP-element group 365: 	 branch_block_stmt_1215/if_stmt_2182_else_link/$entry
      -- CP-element group 365: 	 branch_block_stmt_1215/merge_stmt_2161_PhiAck/$exit
      -- CP-element group 365: 	 branch_block_stmt_1215/merge_stmt_2161_PhiAck/phi_stmt_2162_ack
      -- 
    phi_stmt_2162_ack_6428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2162_ack_0, ack => convolution3D_CP_3583_elements(365)); -- 
    branch_req_5345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(365), ack => if_stmt_2182_branch_req_0); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	227 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	368 
    -- CP-element group 366:  members (2) 
      -- CP-element group 366: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/SplitProtocol/Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/SplitProtocol/Sample/ra
      -- 
    ra_6460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2227_inst_ack_0, ack => convolution3D_CP_3583_elements(366)); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	227 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (2) 
      -- CP-element group 367: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/SplitProtocol/Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/SplitProtocol/Update/ca
      -- 
    ca_6465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2227_inst_ack_1, ack => convolution3D_CP_3583_elements(367)); -- 
    -- CP-element group 368:  join  transition  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	372 
    -- CP-element group 368:  members (5) 
      -- CP-element group 368: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/$exit
      -- CP-element group 368: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/$exit
      -- CP-element group 368: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/$exit
      -- CP-element group 368: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2227/SplitProtocol/$exit
      -- CP-element group 368: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_req
      -- 
    phi_stmt_2221_req_6466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2221_req_6466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(368), ack => phi_stmt_2221_req_1); -- 
    convolution3D_cp_element_group_368: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_368"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(366) & convolution3D_CP_3583_elements(367);
      gj_convolution3D_cp_element_group_368 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	227 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	371 
    -- CP-element group 369:  members (2) 
      -- CP-element group 369: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/SplitProtocol/Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/SplitProtocol/Sample/ra
      -- 
    ra_6483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2220_inst_ack_0, ack => convolution3D_CP_3583_elements(369)); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	227 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (2) 
      -- CP-element group 370: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/SplitProtocol/Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/SplitProtocol/Update/ca
      -- 
    ca_6488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2220_inst_ack_1, ack => convolution3D_CP_3583_elements(370)); -- 
    -- CP-element group 371:  join  transition  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	369 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (5) 
      -- CP-element group 371: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/$exit
      -- CP-element group 371: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/$exit
      -- CP-element group 371: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/$exit
      -- CP-element group 371: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2220/SplitProtocol/$exit
      -- CP-element group 371: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_req
      -- 
    phi_stmt_2214_req_6489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2214_req_6489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(371), ack => phi_stmt_2214_req_1); -- 
    convolution3D_cp_element_group_371: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_371"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(369) & convolution3D_CP_3583_elements(370);
      gj_convolution3D_cp_element_group_371 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(371), clk => clk, reset => reset); --
    end block;
    -- CP-element group 372:  join  transition  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	368 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	376 
    -- CP-element group 372:  members (1) 
      -- CP-element group 372: 	 branch_block_stmt_1215/forx_xbodyx_xi356_forx_xbodyx_xi356_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(368) & convolution3D_CP_3583_elements(371);
      gj_convolution3D_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  transition  output  delay-element  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	221 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (4) 
      -- CP-element group 373: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/$exit
      -- CP-element group 373: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/$exit
      -- CP-element group 373: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_sources/type_cast_2225_konst_delay_trans
      -- CP-element group 373: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2221/phi_stmt_2221_req
      -- 
    phi_stmt_2221_req_6500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2221_req_6500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(373), ack => phi_stmt_2221_req_0); -- 
    -- Element group convolution3D_CP_3583_elements(373) is a control-delay.
    cp_element_373_delay: control_delay_element  generic map(name => " 373_delay", delay_value => 1)  port map(req => convolution3D_CP_3583_elements(221), ack => convolution3D_CP_3583_elements(373), clk => clk, reset =>reset);
    -- CP-element group 374:  transition  output  delay-element  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	221 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (4) 
      -- CP-element group 374: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/$exit
      -- CP-element group 374: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/$exit
      -- CP-element group 374: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_sources/type_cast_2218_konst_delay_trans
      -- CP-element group 374: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/phi_stmt_2214/phi_stmt_2214_req
      -- 
    phi_stmt_2214_req_6508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2214_req_6508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(374), ack => phi_stmt_2214_req_0); -- 
    -- Element group convolution3D_CP_3583_elements(374) is a control-delay.
    cp_element_374_delay: control_delay_element  generic map(name => " 374_delay", delay_value => 1)  port map(req => convolution3D_CP_3583_elements(221), ack => convolution3D_CP_3583_elements(374), clk => clk, reset =>reset);
    -- CP-element group 375:  join  transition  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (1) 
      -- CP-element group 375: 	 branch_block_stmt_1215/forx_xbodyx_xi356x_xpreheader_forx_xbodyx_xi356_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(373) & convolution3D_CP_3583_elements(374);
      gj_convolution3D_cp_element_group_375 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  merge  fork  transition  place  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	372 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376: 	378 
    -- CP-element group 376:  members (2) 
      -- CP-element group 376: 	 branch_block_stmt_1215/merge_stmt_2213_PhiReqMerge
      -- CP-element group 376: 	 branch_block_stmt_1215/merge_stmt_2213_PhiAck/$entry
      -- 
    convolution3D_CP_3583_elements(376) <= OrReduce(convolution3D_CP_3583_elements(372) & convolution3D_CP_3583_elements(375));
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (1) 
      -- CP-element group 377: 	 branch_block_stmt_1215/merge_stmt_2213_PhiAck/phi_stmt_2214_ack
      -- 
    phi_stmt_2214_ack_6513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2214_ack_0, ack => convolution3D_CP_3583_elements(377)); -- 
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	376 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (1) 
      -- CP-element group 378: 	 branch_block_stmt_1215/merge_stmt_2213_PhiAck/phi_stmt_2221_ack
      -- 
    phi_stmt_2221_ack_6514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2221_ack_0, ack => convolution3D_CP_3583_elements(378)); -- 
    -- CP-element group 379:  join  fork  transition  place  output  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	222 
    -- CP-element group 379: 	225 
    -- CP-element group 379:  members (10) 
      -- CP-element group 379: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257__entry__
      -- CP-element group 379: 	 branch_block_stmt_1215/merge_stmt_2213__exit__
      -- CP-element group 379: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/$entry
      -- CP-element group 379: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_sample_start_
      -- CP-element group 379: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/RPIPE_maxpool_input_pipe_2230_Sample/rr
      -- CP-element group 379: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_update_start_
      -- CP-element group 379: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_1215/assign_stmt_2231_to_assign_stmt_2257/type_cast_2234_Update/cr
      -- CP-element group 379: 	 branch_block_stmt_1215/merge_stmt_2213_PhiAck/$exit
      -- 
    rr_5398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(379), ack => RPIPE_maxpool_input_pipe_2230_inst_req_0); -- 
    cr_5417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(379), ack => type_cast_2234_inst_req_1); -- 
    convolution3D_cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_379"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(377) & convolution3D_CP_3583_elements(378);
      gj_convolution3D_cp_element_group_379 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(379), clk => clk, reset => reset); --
    end block;
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	226 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (2) 
      -- CP-element group 380: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/SplitProtocol/Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/SplitProtocol/Sample/ra
      -- 
    ra_6538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2268_inst_ack_0, ack => convolution3D_CP_3583_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	226 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (2) 
      -- CP-element group 381: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/SplitProtocol/Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/SplitProtocol/Update/ca
      -- 
    ca_6543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2268_inst_ack_1, ack => convolution3D_CP_3583_elements(381)); -- 
    -- CP-element group 382:  join  transition  place  output  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (8) 
      -- CP-element group 382: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/$exit
      -- CP-element group 382: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/$exit
      -- CP-element group 382: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/$exit
      -- CP-element group 382: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/$exit
      -- CP-element group 382: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_sources/type_cast_2268/SplitProtocol/$exit
      -- CP-element group 382: 	 branch_block_stmt_1215/forx_xbodyx_xi356_getRemainingElementsx_xexit363_PhiReq/phi_stmt_2265/phi_stmt_2265_req
      -- CP-element group 382: 	 branch_block_stmt_1215/merge_stmt_2264_PhiReqMerge
      -- CP-element group 382: 	 branch_block_stmt_1215/merge_stmt_2264_PhiAck/$entry
      -- 
    phi_stmt_2265_req_6544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2265_req_6544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(382), ack => phi_stmt_2265_req_0); -- 
    convolution3D_cp_element_group_382: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_382"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(380) & convolution3D_CP_3583_elements(381);
      gj_convolution3D_cp_element_group_382 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(382), clk => clk, reset => reset); --
    end block;
    -- CP-element group 383:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	236 
    -- CP-element group 383: 	230 
    -- CP-element group 383: 	231 
    -- CP-element group 383: 	233 
    -- CP-element group 383: 	228 
    -- CP-element group 383: 	229 
    -- CP-element group 383:  members (35) 
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307__entry__
      -- CP-element group 383: 	 branch_block_stmt_1215/merge_stmt_2264__exit__
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_Update/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_final_index_sum_regn_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_Update/cr
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_update_start_
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_final_index_sum_regn_Sample/req
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_update_start_
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_final_index_sum_regn_Update/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_final_index_sum_regn_Update/req
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_complete/req
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/addr_of_2302_complete/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_final_index_sum_regn_update_start
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_scale_1/scale_rename_ack
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_scale_1/scale_rename_req
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_scale_1/$exit
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_scale_1/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_resize_1/index_resize_ack
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_resize_1/index_resize_req
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_resize_1/$exit
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_resize_1/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_computed_1
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Update/word_access_complete/word_0/cr
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Update/word_access_complete/word_0/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Update/word_access_complete/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/ptr_deref_2305_Update/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_scaled_1
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_Sample/rr
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/array_obj_ref_2301_index_resized_1
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/$entry
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_sample_start_
      -- CP-element group 383: 	 branch_block_stmt_1215/assign_stmt_2273_to_assign_stmt_2307/type_cast_2272_update_start_
      -- CP-element group 383: 	 branch_block_stmt_1215/merge_stmt_2264_PhiAck/$exit
      -- CP-element group 383: 	 branch_block_stmt_1215/merge_stmt_2264_PhiAck/phi_stmt_2265_ack
      -- 
    phi_stmt_2265_ack_6549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2265_ack_0, ack => convolution3D_CP_3583_elements(383)); -- 
    cr_5453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(383), ack => type_cast_2272_inst_req_1); -- 
    req_5479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(383), ack => array_obj_ref_2301_index_offset_req_0); -- 
    req_5484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(383), ack => array_obj_ref_2301_index_offset_req_1); -- 
    req_5499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(383), ack => addr_of_2302_final_reg_req_1); -- 
    cr_5549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(383), ack => ptr_deref_2305_store_0_req_1); -- 
    rr_5448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(383), ack => type_cast_2272_inst_req_0); -- 
    -- CP-element group 384:  merge  fork  transition  place  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	216 
    -- CP-element group 384: 	237 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	238 
    -- CP-element group 384: 	239 
    -- CP-element group 384: 	240 
    -- CP-element group 384:  members (16) 
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321__entry__
      -- CP-element group 384: 	 branch_block_stmt_1215/merge_stmt_2309__exit__
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_Sample/req
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_Sample/$entry
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/WPIPE_output_pipe_2313_sample_start_
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_Update/ccr
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_Sample/crr
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_Sample/$entry
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_update_start_
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/call_stmt_2312_sample_start_
      -- CP-element group 384: 	 branch_block_stmt_1215/call_stmt_2312_to_assign_stmt_2321/$entry
      -- CP-element group 384: 	 branch_block_stmt_1215/merge_stmt_2309_PhiReqMerge
      -- CP-element group 384: 	 branch_block_stmt_1215/merge_stmt_2309_PhiAck/$entry
      -- CP-element group 384: 	 branch_block_stmt_1215/merge_stmt_2309_PhiAck/$exit
      -- CP-element group 384: 	 branch_block_stmt_1215/merge_stmt_2309_PhiAck/dummy
      -- 
    req_5575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(384), ack => WPIPE_output_pipe_2313_inst_req_0); -- 
    ccr_5566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(384), ack => call_stmt_2312_call_req_1); -- 
    crr_5561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(384), ack => call_stmt_2312_call_req_0); -- 
    convolution3D_CP_3583_elements(384) <= OrReduce(convolution3D_CP_3583_elements(216) & convolution3D_CP_3583_elements(237));
    -- CP-element group 385:  transition  output  delay-element  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	253 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	389 
    -- CP-element group 385:  members (5) 
      -- CP-element group 385: 	 branch_block_stmt_1215/ifx_xend223_whilex_xbody_PhiReq/$exit
      -- CP-element group 385: 	 branch_block_stmt_1215/ifx_xend223_whilex_xbody_PhiReq/phi_stmt_2359/$exit
      -- CP-element group 385: 	 branch_block_stmt_1215/ifx_xend223_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/$exit
      -- CP-element group 385: 	 branch_block_stmt_1215/ifx_xend223_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2363_konst_delay_trans
      -- CP-element group 385: 	 branch_block_stmt_1215/ifx_xend223_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_req
      -- 
    phi_stmt_2359_req_6571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2359_req_6571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(385), ack => phi_stmt_2359_req_0); -- 
    -- Element group convolution3D_CP_3583_elements(385) is a control-delay.
    cp_element_385_delay: control_delay_element  generic map(name => " 385_delay", delay_value => 1)  port map(req => convolution3D_CP_3583_elements(253), ack => convolution3D_CP_3583_elements(385), clk => clk, reset =>reset);
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	264 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	388 
    -- CP-element group 386:  members (2) 
      -- CP-element group 386: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/SplitProtocol/Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/SplitProtocol/Sample/ra
      -- 
    ra_6591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2365_inst_ack_0, ack => convolution3D_CP_3583_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	264 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (2) 
      -- CP-element group 387: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/SplitProtocol/Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/SplitProtocol/Update/ca
      -- 
    ca_6596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2365_inst_ack_1, ack => convolution3D_CP_3583_elements(387)); -- 
    -- CP-element group 388:  join  transition  output  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	387 
    -- CP-element group 388: 	386 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	389 
    -- CP-element group 388:  members (6) 
      -- CP-element group 388: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 388: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/$exit
      -- CP-element group 388: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/$exit
      -- CP-element group 388: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/$exit
      -- CP-element group 388: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_sources/type_cast_2365/SplitProtocol/$exit
      -- CP-element group 388: 	 branch_block_stmt_1215/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2359/phi_stmt_2359_req
      -- 
    phi_stmt_2359_req_6597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2359_req_6597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(388), ack => phi_stmt_2359_req_1); -- 
    convolution3D_cp_element_group_388: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_388"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3583_elements(387) & convolution3D_CP_3583_elements(386);
      gj_convolution3D_cp_element_group_388 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3583_elements(388), clk => clk, reset => reset); --
    end block;
    -- CP-element group 389:  merge  transition  place  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	388 
    -- CP-element group 389: 	385 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (2) 
      -- CP-element group 389: 	 branch_block_stmt_1215/merge_stmt_2358_PhiAck/$entry
      -- CP-element group 389: 	 branch_block_stmt_1215/merge_stmt_2358_PhiReqMerge
      -- 
    convolution3D_CP_3583_elements(389) <= OrReduce(convolution3D_CP_3583_elements(388) & convolution3D_CP_3583_elements(385));
    -- CP-element group 390:  fork  transition  place  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	254 
    -- CP-element group 390: 	258 
    -- CP-element group 390: 	259 
    -- CP-element group 390: 	260 
    -- CP-element group 390: 	261 
    -- CP-element group 390:  members (20) 
      -- CP-element group 390: 	 branch_block_stmt_1215/merge_stmt_2358__exit__
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401__entry__
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_Sample/req
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_Update/ccr
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/WPIPE_num_out_pipe_2372_sample_start_
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/$entry
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_Sample/crr
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_update_start_
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2390_sample_start_
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_Update/ccr
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_Sample/crr
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_update_start_
      -- CP-element group 390: 	 branch_block_stmt_1215/assign_stmt_2371_to_assign_stmt_2401/call_stmt_2386_sample_start_
      -- CP-element group 390: 	 branch_block_stmt_1215/merge_stmt_2358_PhiAck/phi_stmt_2359_ack
      -- CP-element group 390: 	 branch_block_stmt_1215/merge_stmt_2358_PhiAck/$exit
      -- 
    phi_stmt_2359_ack_6602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2359_ack_0, ack => convolution3D_CP_3583_elements(390)); -- 
    req_5665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(390), ack => WPIPE_num_out_pipe_2372_inst_req_0); -- 
    ccr_5712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(390), ack => call_stmt_2390_call_req_1); -- 
    crr_5707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(390), ack => call_stmt_2390_call_req_0); -- 
    ccr_5698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(390), ack => call_stmt_2386_call_req_1); -- 
    crr_5693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3583_elements(390), ack => call_stmt_2386_call_req_0); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar406_1990_resized : std_logic_vector(13 downto 0);
    signal R_indvar406_1990_scaled : std_logic_vector(13 downto 0);
    signal R_indvar419_1535_resized : std_logic_vector(13 downto 0);
    signal R_indvar419_1535_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1849_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1849_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_2300_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_2300_scaled : std_logic_vector(13 downto 0);
    signal add100_1581 : std_logic_vector(63 downto 0);
    signal add106_1599 : std_logic_vector(63 downto 0);
    signal add112_1617 : std_logic_vector(63 downto 0);
    signal add118_1635 : std_logic_vector(63 downto 0);
    signal add124_1653 : std_logic_vector(63 downto 0);
    signal add130_1671 : std_logic_vector(63 downto 0);
    signal add13_1265 : std_logic_vector(15 downto 0);
    signal add167_2018 : std_logic_vector(63 downto 0);
    signal add173_2036 : std_logic_vector(63 downto 0);
    signal add179_2054 : std_logic_vector(63 downto 0);
    signal add185_2072 : std_logic_vector(63 downto 0);
    signal add191_2090 : std_logic_vector(63 downto 0);
    signal add197_2108 : std_logic_vector(63 downto 0);
    signal add203_2126 : std_logic_vector(63 downto 0);
    signal add23_1290 : std_logic_vector(15 downto 0);
    signal add33_1315 : std_logic_vector(15 downto 0);
    signal add43_1340 : std_logic_vector(15 downto 0);
    signal add53_1365 : std_logic_vector(15 downto 0);
    signal add63_1390 : std_logic_vector(15 downto 0);
    signal add73_1415 : std_logic_vector(15 downto 0);
    signal add94_1563 : std_logic_vector(63 downto 0);
    signal add_1240 : std_logic_vector(31 downto 0);
    signal addx_xi352_2240 : std_logic_vector(63 downto 0);
    signal addx_xi_1789 : std_logic_vector(63 downto 0);
    signal and213_2175 : std_logic_vector(31 downto 0);
    signal and_1720 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1536_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1536_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1536_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1536_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1536_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1536_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1850_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1850_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1850_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1850_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1850_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1850_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1991_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2301_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2301_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2301_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2301_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2301_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2301_root_address : std_logic_vector(13 downto 0);
    signal arrayidx141_1852 : std_logic_vector(31 downto 0);
    signal arrayidx207_1993 : std_logic_vector(31 downto 0);
    signal arrayidx222_2303 : std_logic_vector(31 downto 0);
    signal arrayidx_1538 : std_logic_vector(31 downto 0);
    signal call103_1590 : std_logic_vector(7 downto 0);
    signal call109_1608 : std_logic_vector(7 downto 0);
    signal call115_1626 : std_logic_vector(7 downto 0);
    signal call11_1256 : std_logic_vector(7 downto 0);
    signal call121_1644 : std_logic_vector(7 downto 0);
    signal call127_1662 : std_logic_vector(7 downto 0);
    signal call160_1996 : std_logic_vector(7 downto 0);
    signal call164_2009 : std_logic_vector(7 downto 0);
    signal call16_1268 : std_logic_vector(7 downto 0);
    signal call170_2027 : std_logic_vector(7 downto 0);
    signal call176_2045 : std_logic_vector(7 downto 0);
    signal call182_2063 : std_logic_vector(7 downto 0);
    signal call188_2081 : std_logic_vector(7 downto 0);
    signal call194_2099 : std_logic_vector(7 downto 0);
    signal call200_2117 : std_logic_vector(7 downto 0);
    signal call21_1281 : std_logic_vector(7 downto 0);
    signal call225_2312 : std_logic_vector(63 downto 0);
    signal call266_2417 : std_logic_vector(7 downto 0);
    signal call269_2421 : std_logic_vector(7 downto 0);
    signal call26_1293 : std_logic_vector(7 downto 0);
    signal call271_2424 : std_logic_vector(63 downto 0);
    signal call2_1231 : std_logic_vector(7 downto 0);
    signal call31_1306 : std_logic_vector(7 downto 0);
    signal call36_1318 : std_logic_vector(7 downto 0);
    signal call41_1331 : std_logic_vector(7 downto 0);
    signal call46_1343 : std_logic_vector(7 downto 0);
    signal call51_1356 : std_logic_vector(7 downto 0);
    signal call56_1368 : std_logic_vector(7 downto 0);
    signal call61_1381 : std_logic_vector(7 downto 0);
    signal call66_1393 : std_logic_vector(7 downto 0);
    signal call6_1243 : std_logic_vector(7 downto 0);
    signal call71_1406 : std_logic_vector(7 downto 0);
    signal call87_1541 : std_logic_vector(7 downto 0);
    signal call91_1554 : std_logic_vector(7 downto 0);
    signal call97_1572 : std_logic_vector(7 downto 0);
    signal call_1218 : std_logic_vector(7 downto 0);
    signal callx_xi350_2231 : std_logic_vector(7 downto 0);
    signal callx_xi_1780 : std_logic_vector(7 downto 0);
    signal cmp157365_1891 : std_logic_vector(0 downto 0);
    signal cmp368_1439 : std_logic_vector(0 downto 0);
    signal conv105_1594 : std_logic_vector(63 downto 0);
    signal conv10x_xi358_2273 : std_logic_vector(63 downto 0);
    signal conv10x_xi_1822 : std_logic_vector(63 downto 0);
    signal conv111_1612 : std_logic_vector(63 downto 0);
    signal conv117_1630 : std_logic_vector(63 downto 0);
    signal conv123_1648 : std_logic_vector(63 downto 0);
    signal conv129_1666 : std_logic_vector(63 downto 0);
    signal conv12_1260 : std_logic_vector(15 downto 0);
    signal conv145_1862 : std_logic_vector(31 downto 0);
    signal conv148_1866 : std_logic_vector(31 downto 0);
    signal conv151_1870 : std_logic_vector(31 downto 0);
    signal conv161_2000 : std_logic_vector(63 downto 0);
    signal conv166_2013 : std_logic_vector(63 downto 0);
    signal conv172_2031 : std_logic_vector(63 downto 0);
    signal conv178_2049 : std_logic_vector(63 downto 0);
    signal conv184_2067 : std_logic_vector(63 downto 0);
    signal conv190_2085 : std_logic_vector(63 downto 0);
    signal conv196_2103 : std_logic_vector(63 downto 0);
    signal conv19_1272 : std_logic_vector(15 downto 0);
    signal conv1_1222 : std_logic_vector(31 downto 0);
    signal conv202_2121 : std_logic_vector(63 downto 0);
    signal conv226_2414 : std_logic_vector(63 downto 0);
    signal conv22_1285 : std_logic_vector(15 downto 0);
    signal conv250_2383 : std_logic_vector(63 downto 0);
    signal conv272_2429 : std_logic_vector(63 downto 0);
    signal conv277_2438 : std_logic_vector(31 downto 0);
    signal conv279_2442 : std_logic_vector(31 downto 0);
    signal conv287_2459 : std_logic_vector(7 downto 0);
    signal conv293_2469 : std_logic_vector(7 downto 0);
    signal conv299_2479 : std_logic_vector(7 downto 0);
    signal conv29_1297 : std_logic_vector(15 downto 0);
    signal conv305_2489 : std_logic_vector(7 downto 0);
    signal conv311_2499 : std_logic_vector(7 downto 0);
    signal conv317_2509 : std_logic_vector(7 downto 0);
    signal conv323_2519 : std_logic_vector(7 downto 0);
    signal conv329_2529 : std_logic_vector(7 downto 0);
    signal conv32_1310 : std_logic_vector(15 downto 0);
    signal conv39_1322 : std_logic_vector(15 downto 0);
    signal conv3_1235 : std_logic_vector(31 downto 0);
    signal conv42_1335 : std_logic_vector(15 downto 0);
    signal conv49_1347 : std_logic_vector(15 downto 0);
    signal conv52_1360 : std_logic_vector(15 downto 0);
    signal conv59_1372 : std_logic_vector(15 downto 0);
    signal conv5x_xi351_2235 : std_logic_vector(63 downto 0);
    signal conv5x_xi_1784 : std_logic_vector(63 downto 0);
    signal conv62_1385 : std_logic_vector(15 downto 0);
    signal conv69_1397 : std_logic_vector(15 downto 0);
    signal conv72_1410 : std_logic_vector(15 downto 0);
    signal conv79_1419 : std_logic_vector(31 downto 0);
    signal conv81_1423 : std_logic_vector(31 downto 0);
    signal conv88_1545 : std_logic_vector(63 downto 0);
    signal conv93_1558 : std_logic_vector(63 downto 0);
    signal conv99_1576 : std_logic_vector(63 downto 0);
    signal conv9_1247 : std_logic_vector(15 downto 0);
    signal elementx_x015x_xi349_2221 : std_logic_vector(63 downto 0);
    signal elementx_x015x_xi_1770 : std_logic_vector(63 downto 0);
    signal exitcond12_2401 : std_logic_vector(0 downto 0);
    signal exitcond31_2141 : std_logic_vector(0 downto 0);
    signal exitcond42_1686 : std_logic_vector(0 downto 0);
    signal exitcond6_1806 : std_logic_vector(0 downto 0);
    signal exitcond_2257 : std_logic_vector(0 downto 0);
    signal incx_xi354_2252 : std_logic_vector(7 downto 0);
    signal incx_xi_1801 : std_logic_vector(7 downto 0);
    signal indvar406_1979 : std_logic_vector(63 downto 0);
    signal indvar419_1524 : std_logic_vector(63 downto 0);
    signal indvar_2359 : std_logic_vector(63 downto 0);
    signal indvarx_xnext407_2136 : std_logic_vector(63 downto 0);
    signal indvarx_xnext420_1681 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_2396 : std_logic_vector(63 downto 0);
    signal ix_x0x_xlcssa_1707 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_2162 : std_logic_vector(63 downto 0);
    signal mul146_1875 : std_logic_vector(31 downto 0);
    signal mul149_1880 : std_logic_vector(31 downto 0);
    signal mul152_1885 : std_logic_vector(31 downto 0);
    signal mul249_2371 : std_logic_vector(63 downto 0);
    signal mul280_2447 : std_logic_vector(31 downto 0);
    signal mul283_2452 : std_logic_vector(31 downto 0);
    signal mul82_1433 : std_logic_vector(31 downto 0);
    signal mul_1428 : std_logic_vector(31 downto 0);
    signal mulx_xi360_2285 : std_logic_vector(63 downto 0);
    signal mulx_xi_1834 : std_logic_vector(63 downto 0);
    signal nx_x016x_xi348_2214 : std_logic_vector(7 downto 0);
    signal nx_x016x_xi_1763 : std_logic_vector(7 downto 0);
    signal phitmp372425_2159 : std_logic_vector(63 downto 0);
    signal phitmp426_1704 : std_logic_vector(63 downto 0);
    signal ptr_deref_1673_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1673_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1673_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1673_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1673_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1673_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1854_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1854_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1854_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1854_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1854_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1854_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2128_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2128_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2128_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2128_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2128_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2128_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2305_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2305_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2305_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2305_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2305_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2305_word_offset_0 : std_logic_vector(13 downto 0);
    signal sh_promx_xi361_2291 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1840 : std_logic_vector(63 downto 0);
    signal shl102_1587 : std_logic_vector(63 downto 0);
    signal shl108_1605 : std_logic_vector(63 downto 0);
    signal shl10_1253 : std_logic_vector(15 downto 0);
    signal shl114_1623 : std_logic_vector(63 downto 0);
    signal shl120_1641 : std_logic_vector(63 downto 0);
    signal shl126_1659 : std_logic_vector(63 downto 0);
    signal shl12x_xi362_2296 : std_logic_vector(63 downto 0);
    signal shl12x_xi_1845 : std_logic_vector(63 downto 0);
    signal shl163_2006 : std_logic_vector(63 downto 0);
    signal shl169_2024 : std_logic_vector(63 downto 0);
    signal shl175_2042 : std_logic_vector(63 downto 0);
    signal shl181_2060 : std_logic_vector(63 downto 0);
    signal shl187_2078 : std_logic_vector(63 downto 0);
    signal shl193_2096 : std_logic_vector(63 downto 0);
    signal shl199_2114 : std_logic_vector(63 downto 0);
    signal shl20_1278 : std_logic_vector(15 downto 0);
    signal shl30_1303 : std_logic_vector(15 downto 0);
    signal shl40_1328 : std_logic_vector(15 downto 0);
    signal shl50_1353 : std_logic_vector(15 downto 0);
    signal shl60_1378 : std_logic_vector(15 downto 0);
    signal shl70_1403 : std_logic_vector(15 downto 0);
    signal shl90_1551 : std_logic_vector(63 downto 0);
    signal shl96_1569 : std_logic_vector(63 downto 0);
    signal shl_1228 : std_logic_vector(31 downto 0);
    signal shlx_xi353_2246 : std_logic_vector(63 downto 0);
    signal shlx_xi353x_xlcssa_2265 : std_logic_vector(63 downto 0);
    signal shlx_xi_1795 : std_logic_vector(63 downto 0);
    signal shlx_xix_xlcssa_1814 : std_logic_vector(63 downto 0);
    signal shr290_2465 : std_logic_vector(63 downto 0);
    signal shr296_2475 : std_logic_vector(63 downto 0);
    signal shr302_2485 : std_logic_vector(63 downto 0);
    signal shr308_2495 : std_logic_vector(63 downto 0);
    signal shr314_2505 : std_logic_vector(63 downto 0);
    signal shr320_2515 : std_logic_vector(63 downto 0);
    signal shr326_2525 : std_logic_vector(63 downto 0);
    signal sub_2434 : std_logic_vector(63 downto 0);
    signal subx_xi359_2279 : std_logic_vector(63 downto 0);
    signal subx_xi_1828 : std_logic_vector(63 downto 0);
    signal tmp10_2332 : std_logic_vector(63 downto 0);
    signal tmp11_2338 : std_logic_vector(63 downto 0);
    signal tmp13_2342 : std_logic_vector(63 downto 0);
    signal tmp14_2347 : std_logic_vector(15 downto 0);
    signal tmp15_2351 : std_logic_vector(63 downto 0);
    signal tmp16_2356 : std_logic_vector(63 downto 0);
    signal tmp18_1914 : std_logic_vector(31 downto 0);
    signal tmp19_1918 : std_logic_vector(31 downto 0);
    signal tmp1_1742 : std_logic_vector(31 downto 0);
    signal tmp20_1923 : std_logic_vector(31 downto 0);
    signal tmp21_1927 : std_logic_vector(31 downto 0);
    signal tmp22_1932 : std_logic_vector(31 downto 0);
    signal tmp23_1936 : std_logic_vector(31 downto 0);
    signal tmp24_1941 : std_logic_vector(31 downto 0);
    signal tmp25_1947 : std_logic_vector(31 downto 0);
    signal tmp26_1953 : std_logic_vector(0 downto 0);
    signal tmp28_1966 : std_logic_vector(31 downto 0);
    signal tmp29_1970 : std_logic_vector(63 downto 0);
    signal tmp2_1746 : std_logic_vector(31 downto 0);
    signal tmp30_1976 : std_logic_vector(63 downto 0);
    signal tmp32_1472 : std_logic_vector(31 downto 0);
    signal tmp33_1477 : std_logic_vector(31 downto 0);
    signal tmp34_1481 : std_logic_vector(31 downto 0);
    signal tmp35_1486 : std_logic_vector(31 downto 0);
    signal tmp36_1492 : std_logic_vector(31 downto 0);
    signal tmp37_1498 : std_logic_vector(0 downto 0);
    signal tmp380_2193 : std_logic_vector(7 downto 0);
    signal tmp382_2198 : std_logic_vector(7 downto 0);
    signal tmp384_2203 : std_logic_vector(7 downto 0);
    signal tmp39_1511 : std_logic_vector(31 downto 0);
    signal tmp3_1751 : std_logic_vector(31 downto 0);
    signal tmp404_1904 : std_logic_vector(31 downto 0);
    signal tmp405_1910 : std_logic_vector(0 downto 0);
    signal tmp40_1515 : std_logic_vector(63 downto 0);
    signal tmp413_1451 : std_logic_vector(31 downto 0);
    signal tmp415_1456 : std_logic_vector(31 downto 0);
    signal tmp416_1462 : std_logic_vector(31 downto 0);
    signal tmp417_1468 : std_logic_vector(0 downto 0);
    signal tmp41_1521 : std_logic_vector(63 downto 0);
    signal tmp4_1756 : std_logic_vector(2 downto 0);
    signal tmp5_1760 : std_logic_vector(7 downto 0);
    signal tmp7_2207 : std_logic_vector(2 downto 0);
    signal tmp8_2211 : std_logic_vector(7 downto 0);
    signal tmp9_2328 : std_logic_vector(15 downto 0);
    signal tmp_1737 : std_logic_vector(31 downto 0);
    signal tobool214_2181 : std_logic_vector(0 downto 0);
    signal tobool_1726 : std_logic_vector(0 downto 0);
    signal type_cast_1226_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1251_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1276_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1301_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1326_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1351_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1376_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1401_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1437_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1460_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1466_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1490_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1496_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1503_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1509_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1519_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1528_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1530_wire : std_logic_vector(63 downto 0);
    signal type_cast_1549_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1567_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1585_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1603_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1621_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1639_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1657_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1679_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1698_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1710_wire : std_logic_vector(63 downto 0);
    signal type_cast_1713_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1718_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1724_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1766_wire : std_logic_vector(7 downto 0);
    signal type_cast_1769_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1773_wire : std_logic_vector(63 downto 0);
    signal type_cast_1776_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1793_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1799_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1817_wire : std_logic_vector(63 downto 0);
    signal type_cast_1825_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1832_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1838_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1889_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1902_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1908_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1945_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1951_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1958_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1964_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1974_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1983_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1985_wire : std_logic_vector(63 downto 0);
    signal type_cast_2004_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2022_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2040_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2058_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2076_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2094_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2112_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2134_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2153_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2165_wire : std_logic_vector(63 downto 0);
    signal type_cast_2168_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2173_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2179_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2218_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2220_wire : std_logic_vector(7 downto 0);
    signal type_cast_2225_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2227_wire : std_logic_vector(63 downto 0);
    signal type_cast_2244_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2250_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2268_wire : std_logic_vector(63 downto 0);
    signal type_cast_2276_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2283_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2289_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2326_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2336_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2363_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2365_wire : std_logic_vector(63 downto 0);
    signal type_cast_2381_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2394_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2412_wire : std_logic_vector(63 downto 0);
    signal type_cast_2427_wire : std_logic_vector(63 downto 0);
    signal type_cast_2463_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2473_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2483_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2493_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2503_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2523_wire_constant : std_logic_vector(63 downto 0);
    signal umax27_1960 : std_logic_vector(31 downto 0);
    signal umax38_1505 : std_logic_vector(31 downto 0);
    signal umax418_1700 : std_logic_vector(31 downto 0);
    signal umax_2155 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1536_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1536_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1536_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1536_resized_base_address <= "00000000000000";
    array_obj_ref_1850_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1850_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1850_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1850_resized_base_address <= "00000000000000";
    array_obj_ref_1991_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1991_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1991_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1991_resized_base_address <= "00000000000000";
    array_obj_ref_2301_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2301_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2301_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2301_resized_base_address <= "00000000000000";
    ptr_deref_1673_word_offset_0 <= "00000000000000";
    ptr_deref_1854_word_offset_0 <= "00000000000000";
    ptr_deref_2128_word_offset_0 <= "00000000000000";
    ptr_deref_2305_word_offset_0 <= "00000000000000";
    type_cast_1226_wire_constant <= "00000000000000000000000000001000";
    type_cast_1251_wire_constant <= "0000000000001000";
    type_cast_1276_wire_constant <= "0000000000001000";
    type_cast_1301_wire_constant <= "0000000000001000";
    type_cast_1326_wire_constant <= "0000000000001000";
    type_cast_1351_wire_constant <= "0000000000001000";
    type_cast_1376_wire_constant <= "0000000000001000";
    type_cast_1401_wire_constant <= "0000000000001000";
    type_cast_1437_wire_constant <= "00000000000000000000000000000111";
    type_cast_1460_wire_constant <= "00000000000000000000000000000011";
    type_cast_1466_wire_constant <= "00000000000000000000000000000001";
    type_cast_1490_wire_constant <= "00000000000000000000000000000011";
    type_cast_1496_wire_constant <= "00000000000000000000000000000001";
    type_cast_1503_wire_constant <= "00000000000000000000000000000001";
    type_cast_1509_wire_constant <= "11111111111111111111111111111111";
    type_cast_1519_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1528_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1549_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1567_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1585_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1603_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1621_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1639_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1657_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1679_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1698_wire_constant <= "00000000000000000000000000000001";
    type_cast_1713_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1718_wire_constant <= "00000000000000000000000000000111";
    type_cast_1724_wire_constant <= "00000000000000000000000000000000";
    type_cast_1769_wire_constant <= "00000000";
    type_cast_1776_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1793_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1799_wire_constant <= "00000001";
    type_cast_1825_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    type_cast_1832_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1838_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1889_wire_constant <= "00000000000000000000000000000111";
    type_cast_1902_wire_constant <= "00000000000000000000000000000011";
    type_cast_1908_wire_constant <= "00000000000000000000000000000001";
    type_cast_1945_wire_constant <= "00000000000000000000000000000011";
    type_cast_1951_wire_constant <= "00000000000000000000000000000001";
    type_cast_1958_wire_constant <= "00000000000000000000000000000001";
    type_cast_1964_wire_constant <= "11111111111111111111111111111111";
    type_cast_1974_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1983_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2004_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2022_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2040_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2058_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2076_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2094_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2112_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2134_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2153_wire_constant <= "00000000000000000000000000000001";
    type_cast_2168_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2173_wire_constant <= "00000000000000000000000000000111";
    type_cast_2179_wire_constant <= "00000000000000000000000000000000";
    type_cast_2218_wire_constant <= "00000000";
    type_cast_2225_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2244_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2250_wire_constant <= "00000001";
    type_cast_2276_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    type_cast_2283_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_2289_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2326_wire_constant <= "1111111111111111";
    type_cast_2336_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2363_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2381_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_2394_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2463_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2473_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_2483_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_2493_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2503_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_2513_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2523_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    phi_stmt_1524: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1528_wire_constant & type_cast_1530_wire;
      req <= phi_stmt_1524_req_0 & phi_stmt_1524_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1524",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1524_ack_0,
          idata => idata,
          odata => indvar419_1524,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1524
    phi_stmt_1707: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1710_wire & type_cast_1713_wire_constant;
      req <= phi_stmt_1707_req_0 & phi_stmt_1707_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1707",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1707_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_1707,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1707
    phi_stmt_1763: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1766_wire & type_cast_1769_wire_constant;
      req <= phi_stmt_1763_req_0 & phi_stmt_1763_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1763",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1763_ack_0,
          idata => idata,
          odata => nx_x016x_xi_1763,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1763
    phi_stmt_1770: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1773_wire & type_cast_1776_wire_constant;
      req <= phi_stmt_1770_req_0 & phi_stmt_1770_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1770",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1770_ack_0,
          idata => idata,
          odata => elementx_x015x_xi_1770,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1770
    phi_stmt_1814: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1817_wire;
      req(0) <= phi_stmt_1814_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1814",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1814_ack_0,
          idata => idata,
          odata => shlx_xix_xlcssa_1814,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1814
    phi_stmt_1979: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1983_wire_constant & type_cast_1985_wire;
      req <= phi_stmt_1979_req_0 & phi_stmt_1979_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1979",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1979_ack_0,
          idata => idata,
          odata => indvar406_1979,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1979
    phi_stmt_2162: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2165_wire & type_cast_2168_wire_constant;
      req <= phi_stmt_2162_req_0 & phi_stmt_2162_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2162",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2162_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_2162,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2162
    phi_stmt_2214: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2218_wire_constant & type_cast_2220_wire;
      req <= phi_stmt_2214_req_0 & phi_stmt_2214_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2214",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2214_ack_0,
          idata => idata,
          odata => nx_x016x_xi348_2214,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2214
    phi_stmt_2221: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2225_wire_constant & type_cast_2227_wire;
      req <= phi_stmt_2221_req_0 & phi_stmt_2221_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2221",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2221_ack_0,
          idata => idata,
          odata => elementx_x015x_xi349_2221,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2221
    phi_stmt_2265: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2268_wire;
      req(0) <= phi_stmt_2265_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2265",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2265_ack_0,
          idata => idata,
          odata => shlx_xi353x_xlcssa_2265,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2265
    phi_stmt_2359: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2363_wire_constant & type_cast_2365_wire;
      req <= phi_stmt_2359_req_0 & phi_stmt_2359_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2359",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2359_ack_0,
          idata => idata,
          odata => indvar_2359,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2359
    -- flow-through select operator MUX_1504_inst
    umax38_1505 <= tmp36_1492 when (tmp37_1498(0) /=  '0') else type_cast_1503_wire_constant;
    -- flow-through select operator MUX_1699_inst
    umax418_1700 <= tmp416_1462 when (tmp417_1468(0) /=  '0') else type_cast_1698_wire_constant;
    -- flow-through select operator MUX_1959_inst
    umax27_1960 <= tmp25_1947 when (tmp26_1953(0) /=  '0') else type_cast_1958_wire_constant;
    -- flow-through select operator MUX_2154_inst
    umax_2155 <= tmp404_1904 when (tmp405_1910(0) /=  '0') else type_cast_2153_wire_constant;
    addr_of_1537_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1537_final_reg_req_0;
      addr_of_1537_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1537_final_reg_req_1;
      addr_of_1537_final_reg_ack_1<= rack(0);
      addr_of_1537_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1537_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1536_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1538,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1851_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1851_final_reg_req_0;
      addr_of_1851_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1851_final_reg_req_1;
      addr_of_1851_final_reg_ack_1<= rack(0);
      addr_of_1851_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1851_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1850_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx141_1852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1992_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1992_final_reg_req_0;
      addr_of_1992_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1992_final_reg_req_1;
      addr_of_1992_final_reg_ack_1<= rack(0);
      addr_of_1992_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1992_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1991_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx207_1993,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2302_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2302_final_reg_req_0;
      addr_of_2302_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2302_final_reg_req_1;
      addr_of_2302_final_reg_ack_1<= rack(0);
      addr_of_2302_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2302_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2301_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx222_2303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1221_inst_req_0;
      type_cast_1221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1221_inst_req_1;
      type_cast_1221_inst_ack_1<= rack(0);
      type_cast_1221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1218,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_1222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1234_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1234_inst_req_0;
      type_cast_1234_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1234_inst_req_1;
      type_cast_1234_inst_ack_1<= rack(0);
      type_cast_1234_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1234_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1231,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1235,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1246_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1246_inst_req_0;
      type_cast_1246_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1246_inst_req_1;
      type_cast_1246_inst_ack_1<= rack(0);
      type_cast_1246_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1246_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1243,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_1247,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1259_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1259_inst_req_0;
      type_cast_1259_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1259_inst_req_1;
      type_cast_1259_inst_ack_1<= rack(0);
      type_cast_1259_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1259_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_1256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1260,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1271_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1271_inst_req_0;
      type_cast_1271_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1271_inst_req_1;
      type_cast_1271_inst_ack_1<= rack(0);
      type_cast_1271_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1271_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1268,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_1272,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1284_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1284_inst_req_0;
      type_cast_1284_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1284_inst_req_1;
      type_cast_1284_inst_ack_1<= rack(0);
      type_cast_1284_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1284_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_1281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1296_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1296_inst_req_0;
      type_cast_1296_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1296_inst_req_1;
      type_cast_1296_inst_ack_1<= rack(0);
      type_cast_1296_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1296_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_1293,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1297,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1309_inst_req_0;
      type_cast_1309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1309_inst_req_1;
      type_cast_1309_inst_ack_1<= rack(0);
      type_cast_1309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_1306,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1310,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1321_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1321_inst_req_0;
      type_cast_1321_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1321_inst_req_1;
      type_cast_1321_inst_ack_1<= rack(0);
      type_cast_1321_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1321_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_1318,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1334_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1334_inst_req_0;
      type_cast_1334_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1334_inst_req_1;
      type_cast_1334_inst_ack_1<= rack(0);
      type_cast_1334_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1334_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_1331,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_1335,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1346_inst_req_0;
      type_cast_1346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1346_inst_req_1;
      type_cast_1346_inst_ack_1<= rack(0);
      type_cast_1346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_1343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_1347,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1359_inst_req_0;
      type_cast_1359_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1359_inst_req_1;
      type_cast_1359_inst_ack_1<= rack(0);
      type_cast_1359_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1359_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_1356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_1360,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1371_inst_req_0;
      type_cast_1371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1371_inst_req_1;
      type_cast_1371_inst_ack_1<= rack(0);
      type_cast_1371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_1368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_1372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1384_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1384_inst_req_0;
      type_cast_1384_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1384_inst_req_1;
      type_cast_1384_inst_ack_1<= rack(0);
      type_cast_1384_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1384_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_1381,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_1385,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1396_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1396_inst_req_0;
      type_cast_1396_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1396_inst_req_1;
      type_cast_1396_inst_ack_1<= rack(0);
      type_cast_1396_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1396_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_1393,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1397,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1409_inst_req_0;
      type_cast_1409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1409_inst_req_1;
      type_cast_1409_inst_ack_1<= rack(0);
      type_cast_1409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1409_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_1406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_1410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1418_inst_req_0;
      type_cast_1418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1418_inst_req_1;
      type_cast_1418_inst_ack_1<= rack(0);
      type_cast_1418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1265,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_1419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1422_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1422_inst_req_0;
      type_cast_1422_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1422_inst_req_1;
      type_cast_1422_inst_ack_1<= rack(0);
      type_cast_1422_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1422_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_1423,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1471_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1471_inst_req_0;
      type_cast_1471_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1471_inst_req_1;
      type_cast_1471_inst_ack_1<= rack(0);
      type_cast_1471_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1471_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1265,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp32_1472,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1480_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1480_inst_req_0;
      type_cast_1480_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1480_inst_req_1;
      type_cast_1480_inst_ack_1<= rack(0);
      type_cast_1480_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1480_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp34_1481,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1514_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1514_inst_req_0;
      type_cast_1514_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1514_inst_req_1;
      type_cast_1514_inst_ack_1<= rack(0);
      type_cast_1514_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1514_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp39_1511,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp40_1515,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1530_inst_req_0;
      type_cast_1530_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1530_inst_req_1;
      type_cast_1530_inst_ack_1<= rack(0);
      type_cast_1530_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1530_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext420_1681,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1530_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1544_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1544_inst_req_0;
      type_cast_1544_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1544_inst_req_1;
      type_cast_1544_inst_ack_1<= rack(0);
      type_cast_1544_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1544_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call87_1541,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_1545,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1557_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1557_inst_req_0;
      type_cast_1557_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1557_inst_req_1;
      type_cast_1557_inst_ack_1<= rack(0);
      type_cast_1557_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1557_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call91_1554,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv93_1558,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1575_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1575_inst_req_0;
      type_cast_1575_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1575_inst_req_1;
      type_cast_1575_inst_ack_1<= rack(0);
      type_cast_1575_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1575_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_1572,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_1576,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1593_inst_req_0;
      type_cast_1593_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1593_inst_req_1;
      type_cast_1593_inst_ack_1<= rack(0);
      type_cast_1593_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1593_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call103_1590,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv105_1594,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1611_inst_req_0;
      type_cast_1611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1611_inst_req_1;
      type_cast_1611_inst_ack_1<= rack(0);
      type_cast_1611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call109_1608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv111_1612,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1629_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1629_inst_req_0;
      type_cast_1629_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1629_inst_req_1;
      type_cast_1629_inst_ack_1<= rack(0);
      type_cast_1629_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1629_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_1626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv117_1630,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1647_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1647_inst_req_0;
      type_cast_1647_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1647_inst_req_1;
      type_cast_1647_inst_ack_1<= rack(0);
      type_cast_1647_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1647_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call121_1644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv123_1648,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1665_inst_req_0;
      type_cast_1665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1665_inst_req_1;
      type_cast_1665_inst_ack_1<= rack(0);
      type_cast_1665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1665_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call127_1662,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv129_1666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1703_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1703_inst_req_0;
      type_cast_1703_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1703_inst_req_1;
      type_cast_1703_inst_ack_1<= rack(0);
      type_cast_1703_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1703_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => umax418_1700,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => phitmp426_1704,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1710_inst_req_0;
      type_cast_1710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1710_inst_req_1;
      type_cast_1710_inst_ack_1<= rack(0);
      type_cast_1710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp426_1704,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1710_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1736_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1736_inst_req_0;
      type_cast_1736_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1736_inst_req_1;
      type_cast_1736_inst_ack_1<= rack(0);
      type_cast_1736_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1736_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1265,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp_1737,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1745_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1745_inst_req_0;
      type_cast_1745_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1745_inst_req_1;
      type_cast_1745_inst_ack_1<= rack(0);
      type_cast_1745_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1745_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp2_1746,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1755_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1755_inst_req_0;
      type_cast_1755_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1755_inst_req_1;
      type_cast_1755_inst_ack_1<= rack(0);
      type_cast_1755_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1755_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_1751,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp4_1756,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1759_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1759_inst_req_0;
      type_cast_1759_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1759_inst_req_1;
      type_cast_1759_inst_ack_1<= rack(0);
      type_cast_1759_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1759_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_1756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp5_1760,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1766_inst_req_0;
      type_cast_1766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1766_inst_req_1;
      type_cast_1766_inst_ack_1<= rack(0);
      type_cast_1766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => incx_xi_1801,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1766_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1773_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1773_inst_req_0;
      type_cast_1773_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1773_inst_req_1;
      type_cast_1773_inst_ack_1<= rack(0);
      type_cast_1773_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1773_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shlx_xi_1795,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1773_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1783_inst_req_0;
      type_cast_1783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1783_inst_req_1;
      type_cast_1783_inst_ack_1<= rack(0);
      type_cast_1783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1783_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_1784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1817_inst_req_0;
      type_cast_1817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1817_inst_req_1;
      type_cast_1817_inst_ack_1<= rack(0);
      type_cast_1817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shlx_xi_1795,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1817_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1821_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1821_inst_req_0;
      type_cast_1821_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1821_inst_req_1;
      type_cast_1821_inst_ack_1<= rack(0);
      type_cast_1821_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1821_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul82_1433,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10x_xi_1822,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1861_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1861_inst_req_0;
      type_cast_1861_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1861_inst_req_1;
      type_cast_1861_inst_ack_1<= rack(0);
      type_cast_1861_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1861_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_1415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1862,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1865_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1865_inst_req_0;
      type_cast_1865_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1865_inst_req_1;
      type_cast_1865_inst_ack_1<= rack(0);
      type_cast_1865_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1865_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_1390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv148_1866,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1869_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1869_inst_req_0;
      type_cast_1869_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1869_inst_req_1;
      type_cast_1869_inst_ack_1<= rack(0);
      type_cast_1869_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1869_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv151_1870,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1913_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1913_inst_req_0;
      type_cast_1913_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1913_inst_req_1;
      type_cast_1913_inst_ack_1<= rack(0);
      type_cast_1913_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1913_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp18_1914,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1917_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1917_inst_req_0;
      type_cast_1917_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1917_inst_req_1;
      type_cast_1917_inst_ack_1<= rack(0);
      type_cast_1917_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1917_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1290,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp19_1918,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1926_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1926_inst_req_0;
      type_cast_1926_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1926_inst_req_1;
      type_cast_1926_inst_ack_1<= rack(0);
      type_cast_1926_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1926_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_1390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp21_1927,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1935_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1935_inst_req_0;
      type_cast_1935_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1935_inst_req_1;
      type_cast_1935_inst_ack_1<= rack(0);
      type_cast_1935_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1935_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_1415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp23_1936,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1969_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1969_inst_req_0;
      type_cast_1969_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1969_inst_req_1;
      type_cast_1969_inst_ack_1<= rack(0);
      type_cast_1969_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1969_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp28_1966,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp29_1970,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1985_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1985_inst_req_0;
      type_cast_1985_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1985_inst_req_1;
      type_cast_1985_inst_ack_1<= rack(0);
      type_cast_1985_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1985_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext407_2136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1985_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1999_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1999_inst_req_0;
      type_cast_1999_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1999_inst_req_1;
      type_cast_1999_inst_ack_1<= rack(0);
      type_cast_1999_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1999_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call160_1996,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_2000,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2012_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2012_inst_req_0;
      type_cast_2012_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2012_inst_req_1;
      type_cast_2012_inst_ack_1<= rack(0);
      type_cast_2012_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2012_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_2009,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv166_2013,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2030_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2030_inst_req_0;
      type_cast_2030_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2030_inst_req_1;
      type_cast_2030_inst_ack_1<= rack(0);
      type_cast_2030_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2030_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call170_2027,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv172_2031,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2048_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2048_inst_req_0;
      type_cast_2048_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2048_inst_req_1;
      type_cast_2048_inst_ack_1<= rack(0);
      type_cast_2048_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2048_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call176_2045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv178_2049,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2066_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2066_inst_req_0;
      type_cast_2066_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2066_inst_req_1;
      type_cast_2066_inst_ack_1<= rack(0);
      type_cast_2066_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2066_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call182_2063,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv184_2067,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2084_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2084_inst_req_0;
      type_cast_2084_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2084_inst_req_1;
      type_cast_2084_inst_ack_1<= rack(0);
      type_cast_2084_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2084_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call188_2081,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv190_2085,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2102_inst_req_0;
      type_cast_2102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2102_inst_req_1;
      type_cast_2102_inst_ack_1<= rack(0);
      type_cast_2102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call194_2099,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv196_2103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2120_inst_req_0;
      type_cast_2120_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2120_inst_req_1;
      type_cast_2120_inst_ack_1<= rack(0);
      type_cast_2120_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call200_2117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv202_2121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2158_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2158_inst_req_0;
      type_cast_2158_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2158_inst_req_1;
      type_cast_2158_inst_ack_1<= rack(0);
      type_cast_2158_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2158_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => umax_2155,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => phitmp372425_2159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2165_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2165_inst_req_0;
      type_cast_2165_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2165_inst_req_1;
      type_cast_2165_inst_ack_1<= rack(0);
      type_cast_2165_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2165_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp372425_2159,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2165_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2206_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2206_inst_req_0;
      type_cast_2206_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2206_inst_req_1;
      type_cast_2206_inst_ack_1<= rack(0);
      type_cast_2206_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2206_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp384_2203,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp7_2207,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2210_inst_req_0;
      type_cast_2210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2210_inst_req_1;
      type_cast_2210_inst_ack_1<= rack(0);
      type_cast_2210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp7_2207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp8_2211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2220_inst_req_0;
      type_cast_2220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2220_inst_req_1;
      type_cast_2220_inst_ack_1<= rack(0);
      type_cast_2220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => incx_xi354_2252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2220_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2227_inst_req_0;
      type_cast_2227_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2227_inst_req_1;
      type_cast_2227_inst_ack_1<= rack(0);
      type_cast_2227_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2227_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shlx_xi353_2246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2227_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2234_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2234_inst_req_0;
      type_cast_2234_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2234_inst_req_1;
      type_cast_2234_inst_ack_1<= rack(0);
      type_cast_2234_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2234_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi350_2231,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi351_2235,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2268_inst_req_0;
      type_cast_2268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2268_inst_req_1;
      type_cast_2268_inst_ack_1<= rack(0);
      type_cast_2268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shlx_xi353_2246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2268_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2272_inst_req_0;
      type_cast_2272_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2272_inst_req_1;
      type_cast_2272_inst_ack_1<= rack(0);
      type_cast_2272_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2272_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul152_1885,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10x_xi358_2273,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2331_inst_req_0;
      type_cast_2331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2331_inst_req_1;
      type_cast_2331_inst_ack_1<= rack(0);
      type_cast_2331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp9_2328,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10_2332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2341_inst_req_0;
      type_cast_2341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2341_inst_req_1;
      type_cast_2341_inst_ack_1<= rack(0);
      type_cast_2341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_1390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_2342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2350_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2350_inst_req_0;
      type_cast_2350_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2350_inst_req_1;
      type_cast_2350_inst_ack_1<= rack(0);
      type_cast_2350_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2350_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_2347,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_2351,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2365_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2365_inst_req_0;
      type_cast_2365_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2365_inst_req_1;
      type_cast_2365_inst_ack_1<= rack(0);
      type_cast_2365_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2365_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2365_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2413_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2413_inst_req_0;
      type_cast_2413_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2413_inst_req_1;
      type_cast_2413_inst_ack_1<= rack(0);
      type_cast_2413_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2413_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2412_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv226_2414,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2428_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2428_inst_req_0;
      type_cast_2428_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2428_inst_req_1;
      type_cast_2428_inst_ack_1<= rack(0);
      type_cast_2428_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2428_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2427_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv272_2429,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2437_inst_req_0;
      type_cast_2437_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2437_inst_req_1;
      type_cast_2437_inst_ack_1<= rack(0);
      type_cast_2437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add43_1340,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv277_2438,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2441_inst_req_0;
      type_cast_2441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2441_inst_req_1;
      type_cast_2441_inst_ack_1<= rack(0);
      type_cast_2441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add33_1315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv279_2442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2458_inst_req_0;
      type_cast_2458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2458_inst_req_1;
      type_cast_2458_inst_ack_1<= rack(0);
      type_cast_2458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2458_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_2434,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv287_2459,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2468_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2468_inst_req_0;
      type_cast_2468_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2468_inst_req_1;
      type_cast_2468_inst_ack_1<= rack(0);
      type_cast_2468_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2468_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr290_2465,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv293_2469,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2478_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2478_inst_req_0;
      type_cast_2478_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2478_inst_req_1;
      type_cast_2478_inst_ack_1<= rack(0);
      type_cast_2478_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2478_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr296_2475,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv299_2479,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2488_inst_req_0;
      type_cast_2488_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2488_inst_req_1;
      type_cast_2488_inst_ack_1<= rack(0);
      type_cast_2488_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr302_2485,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_2489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2498_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2498_inst_req_0;
      type_cast_2498_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2498_inst_req_1;
      type_cast_2498_inst_ack_1<= rack(0);
      type_cast_2498_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2498_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr308_2495,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv311_2499,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2508_inst_req_0;
      type_cast_2508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2508_inst_req_1;
      type_cast_2508_inst_ack_1<= rack(0);
      type_cast_2508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr314_2505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv317_2509,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2518_inst_req_0;
      type_cast_2518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2518_inst_req_1;
      type_cast_2518_inst_ack_1<= rack(0);
      type_cast_2518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr320_2515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv323_2519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2528_inst_req_0;
      type_cast_2528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2528_inst_req_1;
      type_cast_2528_inst_ack_1<= rack(0);
      type_cast_2528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr326_2525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv329_2529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1536_index_1_rename
    process(R_indvar419_1535_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar419_1535_resized;
      ov(13 downto 0) := iv;
      R_indvar419_1535_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1536_index_1_resize
    process(indvar419_1524) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar419_1524;
      ov := iv(13 downto 0);
      R_indvar419_1535_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1536_root_address_inst
    process(array_obj_ref_1536_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1536_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1536_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1850_index_1_rename
    process(R_ix_x0x_xlcssa_1849_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1849_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1849_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1850_index_1_resize
    process(ix_x0x_xlcssa_1707) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_1707;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1849_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1850_root_address_inst
    process(array_obj_ref_1850_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1850_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1850_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1991_index_1_rename
    process(R_indvar406_1990_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar406_1990_resized;
      ov(13 downto 0) := iv;
      R_indvar406_1990_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1991_index_1_resize
    process(indvar406_1979) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar406_1979;
      ov := iv(13 downto 0);
      R_indvar406_1990_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1991_root_address_inst
    process(array_obj_ref_1991_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1991_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1991_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2301_index_1_rename
    process(R_ix_x1x_xlcssa_2300_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_2300_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_2300_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2301_index_1_resize
    process(ix_x1x_xlcssa_2162) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_2162;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_2300_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2301_root_address_inst
    process(array_obj_ref_2301_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2301_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2301_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1673_addr_0
    process(ptr_deref_1673_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1673_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1673_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1673_base_resize
    process(arrayidx_1538) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1538;
      ov := iv(13 downto 0);
      ptr_deref_1673_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1673_gather_scatter
    process(add130_1671) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add130_1671;
      ov(63 downto 0) := iv;
      ptr_deref_1673_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1673_root_address_inst
    process(ptr_deref_1673_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1673_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1673_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1854_addr_0
    process(ptr_deref_1854_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1854_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1854_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1854_base_resize
    process(arrayidx141_1852) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx141_1852;
      ov := iv(13 downto 0);
      ptr_deref_1854_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1854_gather_scatter
    process(shl12x_xi_1845) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl12x_xi_1845;
      ov(63 downto 0) := iv;
      ptr_deref_1854_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1854_root_address_inst
    process(ptr_deref_1854_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1854_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1854_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2128_addr_0
    process(ptr_deref_2128_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2128_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2128_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2128_base_resize
    process(arrayidx207_1993) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx207_1993;
      ov := iv(13 downto 0);
      ptr_deref_2128_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2128_gather_scatter
    process(add203_2126) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add203_2126;
      ov(63 downto 0) := iv;
      ptr_deref_2128_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2128_root_address_inst
    process(ptr_deref_2128_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2128_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2128_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2305_addr_0
    process(ptr_deref_2305_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2305_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2305_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2305_base_resize
    process(arrayidx222_2303) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx222_2303;
      ov := iv(13 downto 0);
      ptr_deref_2305_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2305_gather_scatter
    process(shl12x_xi362_2296) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl12x_xi362_2296;
      ov(63 downto 0) := iv;
      ptr_deref_2305_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2305_root_address_inst
    process(ptr_deref_2305_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2305_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2305_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1440_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp368_1439;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1440_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1440_branch_req_0,
          ack0 => if_stmt_1440_branch_ack_0,
          ack1 => if_stmt_1440_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1687_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond42_1686;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1687_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1687_branch_req_0,
          ack0 => if_stmt_1687_branch_ack_0,
          ack1 => if_stmt_1687_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1727_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_1726;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1727_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1727_branch_req_0,
          ack0 => if_stmt_1727_branch_ack_0,
          ack1 => if_stmt_1727_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1807_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond6_1806;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1807_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1807_branch_req_0,
          ack0 => if_stmt_1807_branch_ack_0,
          ack1 => if_stmt_1807_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1892_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp157365_1891;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1892_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1892_branch_req_0,
          ack0 => if_stmt_1892_branch_ack_0,
          ack1 => if_stmt_1892_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2142_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond31_2141;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2142_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2142_branch_req_0,
          ack0 => if_stmt_2142_branch_ack_0,
          ack1 => if_stmt_2142_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2182_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool214_2181;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2182_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2182_branch_req_0,
          ack0 => if_stmt_2182_branch_ack_0,
          ack1 => if_stmt_2182_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2258_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_2257;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2258_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2258_branch_req_0,
          ack0 => if_stmt_2258_branch_ack_0,
          ack1 => if_stmt_2258_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2402_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond12_2401;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2402_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2402_branch_req_0,
          ack0 => if_stmt_2402_branch_ack_0,
          ack1 => if_stmt_2402_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2327_inst
    process(add53_1365) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_1365, type_cast_2326_wire_constant, tmp_var);
      tmp9_2328 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1510_inst
    process(umax38_1505) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(umax38_1505, type_cast_1509_wire_constant, tmp_var);
      tmp39_1511 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1965_inst
    process(umax27_1960) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(umax27_1960, type_cast_1964_wire_constant, tmp_var);
      tmp28_1966 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1520_inst
    process(tmp40_1515) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp40_1515, type_cast_1519_wire_constant, tmp_var);
      tmp41_1521 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1680_inst
    process(indvar419_1524) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar419_1524, type_cast_1679_wire_constant, tmp_var);
      indvarx_xnext420_1681 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1975_inst
    process(tmp29_1970) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp29_1970, type_cast_1974_wire_constant, tmp_var);
      tmp30_1976 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2135_inst
    process(indvar406_1979) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar406_1979, type_cast_2134_wire_constant, tmp_var);
      indvarx_xnext407_2136 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2337_inst
    process(tmp10_2332) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp10_2332, type_cast_2336_wire_constant, tmp_var);
      tmp11_2338 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2395_inst
    process(indvar_2359) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2359, type_cast_2394_wire_constant, tmp_var);
      indvarx_xnext_2396 <= tmp_var; --
    end process;
    -- binary operator ADD_u8_u8_1800_inst
    process(nx_x016x_xi_1763) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x016x_xi_1763, type_cast_1799_wire_constant, tmp_var);
      incx_xi_1801 <= tmp_var; --
    end process;
    -- binary operator ADD_u8_u8_2251_inst
    process(nx_x016x_xi348_2214) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x016x_xi348_2214, type_cast_2250_wire_constant, tmp_var);
      incx_xi354_2252 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1719_inst
    process(mul82_1433) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul82_1433, type_cast_1718_wire_constant, tmp_var);
      and_1720 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2174_inst
    process(mul152_1885) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul152_1885, type_cast_2173_wire_constant, tmp_var);
      and213_2175 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1839_inst
    process(mulx_xi_1834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mulx_xi_1834, type_cast_1838_wire_constant, tmp_var);
      sh_promx_xi_1840 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2290_inst
    process(mulx_xi360_2285) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mulx_xi360_2285, type_cast_2289_wire_constant, tmp_var);
      sh_promx_xi361_2291 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2382_inst
    process(mul249_2371) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul249_2371, type_cast_2381_wire_constant, tmp_var);
      conv250_2383 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1725_inst
    process(and_1720) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_1720, type_cast_1724_wire_constant, tmp_var);
      tobool_1726 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2180_inst
    process(and213_2175) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and213_2175, type_cast_2179_wire_constant, tmp_var);
      tobool214_2181 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1685_inst
    process(indvarx_xnext420_1681, tmp41_1521) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext420_1681, tmp41_1521, tmp_var);
      exitcond42_1686 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2140_inst
    process(indvarx_xnext407_2136, tmp30_1976) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext407_2136, tmp30_1976, tmp_var);
      exitcond31_2141 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2400_inst
    process(indvarx_xnext_2396, tmp11_2338) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_2396, tmp11_2338, tmp_var);
      exitcond12_2401 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1805_inst
    process(incx_xi_1801, tmp5_1760) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(incx_xi_1801, tmp5_1760, tmp_var);
      exitcond6_1806 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_2256_inst
    process(incx_xi354_2252, tmp8_2211) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(incx_xi354_2252, tmp8_2211, tmp_var);
      exitcond_2257 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1461_inst
    process(tmp415_1456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp415_1456, type_cast_1460_wire_constant, tmp_var);
      tmp416_1462 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1491_inst
    process(tmp35_1486) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp35_1486, type_cast_1490_wire_constant, tmp_var);
      tmp36_1492 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1903_inst
    process(mul152_1885) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul152_1885, type_cast_1902_wire_constant, tmp_var);
      tmp404_1904 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1946_inst
    process(tmp24_1941) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp24_1941, type_cast_1945_wire_constant, tmp_var);
      tmp25_1947 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2464_inst
    process(sub_2434) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2434, type_cast_2463_wire_constant, tmp_var);
      shr290_2465 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2474_inst
    process(sub_2434) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2434, type_cast_2473_wire_constant, tmp_var);
      shr296_2475 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2484_inst
    process(sub_2434) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2434, type_cast_2483_wire_constant, tmp_var);
      shr302_2485 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2494_inst
    process(sub_2434) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2434, type_cast_2493_wire_constant, tmp_var);
      shr308_2495 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2504_inst
    process(sub_2434) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2434, type_cast_2503_wire_constant, tmp_var);
      shr314_2505 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2514_inst
    process(sub_2434) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2434, type_cast_2513_wire_constant, tmp_var);
      shr320_2515 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2524_inst
    process(sub_2434) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2434, type_cast_2523_wire_constant, tmp_var);
      shr326_2525 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2346_inst
    process(add73_1415, add23_1290) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1415, add23_1290, tmp_var);
      tmp14_2347 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1427_inst
    process(conv79_1419, add_1240) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_1419, add_1240, tmp_var);
      mul_1428 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1432_inst
    process(mul_1428, conv81_1423) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1428, conv81_1423, tmp_var);
      mul82_1433 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1450_inst
    process(add_1240, conv79_1419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1240, conv79_1419, tmp_var);
      tmp413_1451 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1455_inst
    process(tmp413_1451, conv81_1423) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp413_1451, conv81_1423, tmp_var);
      tmp415_1456 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1476_inst
    process(add_1240, tmp32_1472) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1240, tmp32_1472, tmp_var);
      tmp33_1477 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1485_inst
    process(tmp33_1477, tmp34_1481) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp33_1477, tmp34_1481, tmp_var);
      tmp35_1486 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1741_inst
    process(add_1240, tmp_1737) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1240, tmp_1737, tmp_var);
      tmp1_1742 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1750_inst
    process(tmp1_1742, tmp2_1746) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_1742, tmp2_1746, tmp_var);
      tmp3_1751 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1874_inst
    process(conv151_1870, conv81_1423) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv151_1870, conv81_1423, tmp_var);
      mul146_1875 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1879_inst
    process(mul146_1875, conv148_1866) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul146_1875, conv148_1866, tmp_var);
      mul149_1880 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1884_inst
    process(mul149_1880, conv145_1862) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul149_1880, conv145_1862, tmp_var);
      mul152_1885 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1922_inst
    process(tmp18_1914, tmp19_1918) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp18_1914, tmp19_1918, tmp_var);
      tmp20_1923 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1931_inst
    process(tmp20_1923, tmp21_1927) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp20_1923, tmp21_1927, tmp_var);
      tmp22_1932 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1940_inst
    process(tmp22_1932, tmp23_1936) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp22_1932, tmp23_1936, tmp_var);
      tmp24_1941 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2446_inst
    process(conv277_2438, conv279_2442) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv277_2438, conv279_2442, tmp_var);
      mul280_2447 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2451_inst
    process(mul280_2447, conv151_1870) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul280_2447, conv151_1870, tmp_var);
      mul283_2452 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2355_inst
    process(tmp13_2342, tmp15_2351) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_2342, tmp15_2351, tmp_var);
      tmp16_2356 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2370_inst
    process(tmp16_2356, indvar_2359) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_2356, indvar_2359, tmp_var);
      mul249_2371 <= tmp_var; --
    end process;
    -- binary operator MUL_u8_u8_2192_inst
    process(call51_1356, call21_1281) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(call51_1356, call21_1281, tmp_var);
      tmp380_2193 <= tmp_var; --
    end process;
    -- binary operator MUL_u8_u8_2197_inst
    process(tmp380_2193, call61_1381) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp380_2193, call61_1381, tmp_var);
      tmp382_2198 <= tmp_var; --
    end process;
    -- binary operator MUL_u8_u8_2202_inst
    process(tmp382_2198, call71_1406) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp382_2198, call71_1406, tmp_var);
      tmp384_2203 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1264_inst
    process(shl10_1253, conv12_1260) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_1253, conv12_1260, tmp_var);
      add13_1265 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1289_inst
    process(shl20_1278, conv22_1285) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_1278, conv22_1285, tmp_var);
      add23_1290 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1314_inst
    process(shl30_1303, conv32_1310) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_1303, conv32_1310, tmp_var);
      add33_1315 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1339_inst
    process(shl40_1328, conv42_1335) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_1328, conv42_1335, tmp_var);
      add43_1340 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1364_inst
    process(shl50_1353, conv52_1360) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_1353, conv52_1360, tmp_var);
      add53_1365 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1389_inst
    process(shl60_1378, conv62_1385) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_1378, conv62_1385, tmp_var);
      add63_1390 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1414_inst
    process(shl70_1403, conv72_1410) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_1403, conv72_1410, tmp_var);
      add73_1415 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1239_inst
    process(shl_1228, conv3_1235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1228, conv3_1235, tmp_var);
      add_1240 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1562_inst
    process(shl90_1551, conv93_1558) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl90_1551, conv93_1558, tmp_var);
      add94_1563 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1580_inst
    process(shl96_1569, conv99_1576) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_1569, conv99_1576, tmp_var);
      add100_1581 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1598_inst
    process(shl102_1587, conv105_1594) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl102_1587, conv105_1594, tmp_var);
      add106_1599 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1616_inst
    process(shl108_1605, conv111_1612) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl108_1605, conv111_1612, tmp_var);
      add112_1617 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1634_inst
    process(shl114_1623, conv117_1630) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_1623, conv117_1630, tmp_var);
      add118_1635 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1652_inst
    process(shl120_1641, conv123_1648) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl120_1641, conv123_1648, tmp_var);
      add124_1653 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1670_inst
    process(shl126_1659, conv129_1666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl126_1659, conv129_1666, tmp_var);
      add130_1671 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1788_inst
    process(conv5x_xi_1784, elementx_x015x_xi_1770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_1784, elementx_x015x_xi_1770, tmp_var);
      addx_xi_1789 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2017_inst
    process(shl163_2006, conv166_2013) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl163_2006, conv166_2013, tmp_var);
      add167_2018 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2035_inst
    process(shl169_2024, conv172_2031) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl169_2024, conv172_2031, tmp_var);
      add173_2036 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2053_inst
    process(shl175_2042, conv178_2049) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl175_2042, conv178_2049, tmp_var);
      add179_2054 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2071_inst
    process(shl181_2060, conv184_2067) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl181_2060, conv184_2067, tmp_var);
      add185_2072 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2089_inst
    process(shl187_2078, conv190_2085) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl187_2078, conv190_2085, tmp_var);
      add191_2090 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2107_inst
    process(shl193_2096, conv196_2103) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl193_2096, conv196_2103, tmp_var);
      add197_2108 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2125_inst
    process(shl199_2114, conv202_2121) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl199_2114, conv202_2121, tmp_var);
      add203_2126 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2239_inst
    process(conv5x_xi351_2235, elementx_x015x_xi349_2221) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi351_2235, elementx_x015x_xi349_2221, tmp_var);
      addx_xi352_2240 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1252_inst
    process(conv9_1247) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_1247, type_cast_1251_wire_constant, tmp_var);
      shl10_1253 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1277_inst
    process(conv19_1272) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_1272, type_cast_1276_wire_constant, tmp_var);
      shl20_1278 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1302_inst
    process(conv29_1297) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_1297, type_cast_1301_wire_constant, tmp_var);
      shl30_1303 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1327_inst
    process(conv39_1322) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_1322, type_cast_1326_wire_constant, tmp_var);
      shl40_1328 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1352_inst
    process(conv49_1347) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_1347, type_cast_1351_wire_constant, tmp_var);
      shl50_1353 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1377_inst
    process(conv59_1372) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_1372, type_cast_1376_wire_constant, tmp_var);
      shl60_1378 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1402_inst
    process(conv69_1397) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_1397, type_cast_1401_wire_constant, tmp_var);
      shl70_1403 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1227_inst
    process(conv1_1222) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_1222, type_cast_1226_wire_constant, tmp_var);
      shl_1228 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1550_inst
    process(conv88_1545) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv88_1545, type_cast_1549_wire_constant, tmp_var);
      shl90_1551 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1568_inst
    process(add94_1563) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add94_1563, type_cast_1567_wire_constant, tmp_var);
      shl96_1569 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1586_inst
    process(add100_1581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add100_1581, type_cast_1585_wire_constant, tmp_var);
      shl102_1587 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1604_inst
    process(add106_1599) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add106_1599, type_cast_1603_wire_constant, tmp_var);
      shl108_1605 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1622_inst
    process(add112_1617) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add112_1617, type_cast_1621_wire_constant, tmp_var);
      shl114_1623 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1640_inst
    process(add118_1635) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add118_1635, type_cast_1639_wire_constant, tmp_var);
      shl120_1641 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1658_inst
    process(add124_1653) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add124_1653, type_cast_1657_wire_constant, tmp_var);
      shl126_1659 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1794_inst
    process(addx_xi_1789) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1789, type_cast_1793_wire_constant, tmp_var);
      shlx_xi_1795 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1833_inst
    process(subx_xi_1828) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(subx_xi_1828, type_cast_1832_wire_constant, tmp_var);
      mulx_xi_1834 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1844_inst
    process(shlx_xix_xlcssa_1814, sh_promx_xi_1840) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shlx_xix_xlcssa_1814, sh_promx_xi_1840, tmp_var);
      shl12x_xi_1845 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2005_inst
    process(conv161_2000) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv161_2000, type_cast_2004_wire_constant, tmp_var);
      shl163_2006 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2023_inst
    process(add167_2018) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add167_2018, type_cast_2022_wire_constant, tmp_var);
      shl169_2024 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2041_inst
    process(add173_2036) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add173_2036, type_cast_2040_wire_constant, tmp_var);
      shl175_2042 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2059_inst
    process(add179_2054) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add179_2054, type_cast_2058_wire_constant, tmp_var);
      shl181_2060 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2077_inst
    process(add185_2072) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add185_2072, type_cast_2076_wire_constant, tmp_var);
      shl187_2078 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2095_inst
    process(add191_2090) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add191_2090, type_cast_2094_wire_constant, tmp_var);
      shl193_2096 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2113_inst
    process(add197_2108) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add197_2108, type_cast_2112_wire_constant, tmp_var);
      shl199_2114 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2245_inst
    process(addx_xi352_2240) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi352_2240, type_cast_2244_wire_constant, tmp_var);
      shlx_xi353_2246 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2284_inst
    process(subx_xi359_2279) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(subx_xi359_2279, type_cast_2283_wire_constant, tmp_var);
      mulx_xi360_2285 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2295_inst
    process(shlx_xi353x_xlcssa_2265, sh_promx_xi361_2291) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shlx_xi353x_xlcssa_2265, sh_promx_xi361_2291, tmp_var);
      shl12x_xi362_2296 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1827_inst
    process(type_cast_1825_wire_constant, conv10x_xi_1822) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(type_cast_1825_wire_constant, conv10x_xi_1822, tmp_var);
      subx_xi_1828 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_2278_inst
    process(type_cast_2276_wire_constant, conv10x_xi358_2273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(type_cast_2276_wire_constant, conv10x_xi358_2273, tmp_var);
      subx_xi359_2279 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_2433_inst
    process(conv272_2429, conv226_2414) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv272_2429, conv226_2414, tmp_var);
      sub_2434 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1438_inst
    process(mul82_1433) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_1433, type_cast_1437_wire_constant, tmp_var);
      cmp368_1439 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1467_inst
    process(tmp416_1462) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp416_1462, type_cast_1466_wire_constant, tmp_var);
      tmp417_1468 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1497_inst
    process(tmp36_1492) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp36_1492, type_cast_1496_wire_constant, tmp_var);
      tmp37_1498 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1890_inst
    process(mul152_1885) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul152_1885, type_cast_1889_wire_constant, tmp_var);
      cmp157365_1891 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1909_inst
    process(tmp404_1904) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp404_1904, type_cast_1908_wire_constant, tmp_var);
      tmp405_1910 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1952_inst
    process(tmp25_1947) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp25_1947, type_cast_1951_wire_constant, tmp_var);
      tmp26_1953 <= tmp_var; --
    end process;
    -- shared split operator group (117) : array_obj_ref_1536_index_offset 
    ApIntAdd_group_117: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar419_1535_scaled;
      array_obj_ref_1536_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1536_index_offset_req_0;
      array_obj_ref_1536_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1536_index_offset_req_1;
      array_obj_ref_1536_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_117_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_117_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- shared split operator group (118) : array_obj_ref_1850_index_offset 
    ApIntAdd_group_118: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1849_scaled;
      array_obj_ref_1850_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1850_index_offset_req_0;
      array_obj_ref_1850_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1850_index_offset_req_1;
      array_obj_ref_1850_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_118_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_118_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- shared split operator group (119) : array_obj_ref_1991_index_offset 
    ApIntAdd_group_119: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar406_1990_scaled;
      array_obj_ref_1991_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1991_index_offset_req_0;
      array_obj_ref_1991_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1991_index_offset_req_1;
      array_obj_ref_1991_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_119_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_119_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_119",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 119
    -- shared split operator group (120) : array_obj_ref_2301_index_offset 
    ApIntAdd_group_120: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_2300_scaled;
      array_obj_ref_2301_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2301_index_offset_req_0;
      array_obj_ref_2301_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2301_index_offset_req_1;
      array_obj_ref_2301_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_120_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_120_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_120",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 120
    -- unary operator type_cast_2412_inst
    process(call225_2312) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call225_2312, tmp_var);
      type_cast_2412_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2427_inst
    process(call271_2424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call271_2424, tmp_var);
      type_cast_2427_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1854_store_0 ptr_deref_1673_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1854_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1673_store_0_req_0;
      ptr_deref_1854_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1673_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1854_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1673_store_0_req_1;
      ptr_deref_1854_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1673_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1854_word_address_0 & ptr_deref_1673_word_address_0;
      data_in <= ptr_deref_1854_data_0 & ptr_deref_1673_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_2128_store_0 ptr_deref_2305_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2128_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2305_store_0_req_0;
      ptr_deref_2128_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2305_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2128_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2305_store_0_req_1;
      ptr_deref_2128_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2305_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2128_word_address_0 & ptr_deref_2305_word_address_0;
      data_in <= ptr_deref_2128_data_0 & ptr_deref_2305_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_input_done_pipe_2416_inst RPIPE_input_done_pipe_2420_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_input_done_pipe_2416_inst_req_0;
      reqL_unguarded(0) <= RPIPE_input_done_pipe_2420_inst_req_0;
      RPIPE_input_done_pipe_2416_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_input_done_pipe_2420_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_input_done_pipe_2416_inst_req_1;
      reqR_unguarded(0) <= RPIPE_input_done_pipe_2420_inst_req_1;
      RPIPE_input_done_pipe_2416_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_input_done_pipe_2420_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      call266_2417 <= data_out(15 downto 8);
      call269_2421 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_maxpool_input_pipe_1995_inst RPIPE_maxpool_input_pipe_2080_inst RPIPE_maxpool_input_pipe_1589_inst RPIPE_maxpool_input_pipe_1625_inst RPIPE_maxpool_input_pipe_2116_inst RPIPE_maxpool_input_pipe_2008_inst RPIPE_maxpool_input_pipe_1643_inst RPIPE_maxpool_input_pipe_1571_inst RPIPE_maxpool_input_pipe_2026_inst RPIPE_maxpool_input_pipe_1661_inst RPIPE_maxpool_input_pipe_1553_inst RPIPE_maxpool_input_pipe_1540_inst RPIPE_maxpool_input_pipe_2044_inst RPIPE_maxpool_input_pipe_2098_inst RPIPE_maxpool_input_pipe_1607_inst RPIPE_maxpool_input_pipe_1779_inst RPIPE_maxpool_input_pipe_2062_inst RPIPE_maxpool_input_pipe_2230_inst RPIPE_maxpool_input_pipe_1217_inst RPIPE_maxpool_input_pipe_1230_inst RPIPE_maxpool_input_pipe_1242_inst RPIPE_maxpool_input_pipe_1255_inst RPIPE_maxpool_input_pipe_1267_inst RPIPE_maxpool_input_pipe_1280_inst RPIPE_maxpool_input_pipe_1292_inst RPIPE_maxpool_input_pipe_1305_inst RPIPE_maxpool_input_pipe_1317_inst RPIPE_maxpool_input_pipe_1330_inst RPIPE_maxpool_input_pipe_1342_inst RPIPE_maxpool_input_pipe_1355_inst RPIPE_maxpool_input_pipe_1367_inst RPIPE_maxpool_input_pipe_1380_inst RPIPE_maxpool_input_pipe_1392_inst RPIPE_maxpool_input_pipe_1405_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_1995_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_2080_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_1589_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_1625_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_2116_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_2008_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_1643_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_1571_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_2026_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_1661_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_1553_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_1540_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_2044_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_2098_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_1607_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_1779_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_2062_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_2230_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_1217_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_1230_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_1242_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_1255_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_1267_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_1280_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_1292_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_1305_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_1317_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_1330_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_1342_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_1355_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_1367_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_1380_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1392_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1405_inst_req_0;
      RPIPE_maxpool_input_pipe_1995_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_2080_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_1589_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_1625_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_2116_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_2008_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_1643_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_1571_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_2026_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_1661_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_1553_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_1540_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_2044_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_2098_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_1607_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_1779_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_2062_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_2230_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_1217_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_1230_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_1242_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_1255_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_1267_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_1280_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_1292_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_1305_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_1317_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_1330_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_1342_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_1355_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_1367_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_1380_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1392_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1405_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_1995_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_2080_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_1589_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_1625_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_2116_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_2008_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_1643_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_1571_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_2026_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_1661_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_1553_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_1540_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_2044_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_2098_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_1607_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_1779_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_2062_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_2230_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_1217_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_1230_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_1242_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_1255_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_1267_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_1280_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_1292_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_1305_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_1317_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_1330_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_1342_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_1355_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_1367_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_1380_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1392_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1405_inst_req_1;
      RPIPE_maxpool_input_pipe_1995_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_2080_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_1589_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_1625_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_2116_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_2008_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_1643_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_1571_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_2026_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_1661_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_1553_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_1540_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_2044_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_2098_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_1607_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_1779_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_2062_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_2230_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_1217_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_1230_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_1242_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_1255_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_1267_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_1280_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_1292_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_1305_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_1317_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_1330_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_1342_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_1355_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_1367_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_1380_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1392_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1405_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call160_1996 <= data_out(271 downto 264);
      call188_2081 <= data_out(263 downto 256);
      call103_1590 <= data_out(255 downto 248);
      call115_1626 <= data_out(247 downto 240);
      call200_2117 <= data_out(239 downto 232);
      call164_2009 <= data_out(231 downto 224);
      call121_1644 <= data_out(223 downto 216);
      call97_1572 <= data_out(215 downto 208);
      call170_2027 <= data_out(207 downto 200);
      call127_1662 <= data_out(199 downto 192);
      call91_1554 <= data_out(191 downto 184);
      call87_1541 <= data_out(183 downto 176);
      call176_2045 <= data_out(175 downto 168);
      call194_2099 <= data_out(167 downto 160);
      call109_1608 <= data_out(159 downto 152);
      callx_xi_1780 <= data_out(151 downto 144);
      call182_2063 <= data_out(143 downto 136);
      callx_xi350_2231 <= data_out(135 downto 128);
      call_1218 <= data_out(127 downto 120);
      call2_1231 <= data_out(119 downto 112);
      call6_1243 <= data_out(111 downto 104);
      call11_1256 <= data_out(103 downto 96);
      call16_1268 <= data_out(95 downto 88);
      call21_1281 <= data_out(87 downto 80);
      call26_1293 <= data_out(79 downto 72);
      call31_1306 <= data_out(71 downto 64);
      call36_1318 <= data_out(63 downto 56);
      call41_1331 <= data_out(55 downto 48);
      call46_1343 <= data_out(47 downto 40);
      call51_1356 <= data_out(39 downto 32);
      call56_1368 <= data_out(31 downto 24);
      call61_1381 <= data_out(23 downto 16);
      call66_1393 <= data_out(15 downto 8);
      call71_1406 <= data_out(7 downto 0);
      maxpool_input_pipe_read_1_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_1_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_1: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_1", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_2530_inst WPIPE_maxpool_output_pipe_2533_inst WPIPE_maxpool_output_pipe_2536_inst WPIPE_maxpool_output_pipe_2539_inst WPIPE_maxpool_output_pipe_2542_inst WPIPE_maxpool_output_pipe_2545_inst WPIPE_maxpool_output_pipe_2548_inst WPIPE_maxpool_output_pipe_2551_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_2530_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_2533_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_2536_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_2539_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_2542_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_2545_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_2548_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2551_inst_req_0;
      WPIPE_maxpool_output_pipe_2530_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_2533_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_2536_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_2539_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_2542_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_2545_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_2548_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2551_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_2530_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_2533_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_2536_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_2539_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_2542_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_2545_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_2548_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2551_inst_req_1;
      WPIPE_maxpool_output_pipe_2530_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_2533_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_2536_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_2539_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_2542_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_2545_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_2548_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2551_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv329_2529 & conv323_2519 & conv317_2509 & conv311_2499 & conv305_2489 & conv299_2479 & conv293_2469 & conv287_2459;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_num_out_pipe_2372_inst WPIPE_num_out_pipe_2375_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_num_out_pipe_2372_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_2375_inst_req_0;
      WPIPE_num_out_pipe_2372_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_num_out_pipe_2375_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_num_out_pipe_2372_inst_req_1;
      update_req_unguarded(0) <= WPIPE_num_out_pipe_2375_inst_req_1;
      WPIPE_num_out_pipe_2372_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_num_out_pipe_2375_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= add33_1315 & add43_1340;
      num_out_pipe_write_1_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_output_pipe_2313_inst WPIPE_output_pipe_2316_inst WPIPE_output_pipe_2319_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal sample_req, sample_ack : BooleanArray( 2 downto 0);
      signal update_req, update_ack : BooleanArray( 2 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 2 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      sample_req_unguarded(2) <= WPIPE_output_pipe_2313_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_output_pipe_2316_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_output_pipe_2319_inst_req_0;
      WPIPE_output_pipe_2313_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_output_pipe_2316_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_output_pipe_2319_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(2) <= WPIPE_output_pipe_2313_inst_req_1;
      update_req_unguarded(1) <= WPIPE_output_pipe_2316_inst_req_1;
      update_req_unguarded(0) <= WPIPE_output_pipe_2319_inst_req_1;
      WPIPE_output_pipe_2313_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_output_pipe_2316_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_output_pipe_2319_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      data_in <= add33_1315 & add43_1340 & add53_1365;
      output_pipe_write_2_gI: SplitGuardInterface generic map(name => "output_pipe_write_2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "output_pipe", data_width => 16, num_reqs => 3, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => output_pipe_pipe_write_req(0),
          oack => output_pipe_pipe_write_ack(0),
          odata => output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_2312_call call_stmt_2424_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_2312_call_req_0;
      reqL_unguarded(0) <= call_stmt_2424_call_req_0;
      call_stmt_2312_call_ack_0 <= ackL_unguarded(1);
      call_stmt_2424_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_2312_call_req_1;
      reqR_unguarded(0) <= call_stmt_2424_call_req_1;
      call_stmt_2312_call_ack_1 <= ackR_unguarded(1);
      call_stmt_2424_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call225_2312 <= data_out(127 downto 64);
      call271_2424 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2386_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2386_call_req_0;
      call_stmt_2386_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2386_call_req_1;
      call_stmt_2386_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv250_2383 & add23_1290;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(79 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_2390_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2390_call_req_0;
      call_stmt_2390_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2390_call_req_1;
      call_stmt_2390_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= add33_1315 & add23_1290 & add13_1265;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 48,
        owidth => 48,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(47 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_2454_call 
    sendB_call_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2454_call_req_0;
      call_stmt_2454_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2454_call_req_1;
      call_stmt_2454_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendB_call_group_3_gI: SplitGuardInterface generic map(name => "sendB_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul283_2452;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendB_call_reqs(0),
          ackR => sendB_call_acks(0),
          dataR => sendB_call_data(31 downto 0),
          tagR => sendB_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendB_return_acks(0), -- cross-over
          ackL => sendB_return_reqs(0), -- cross-over
          tagL => sendB_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_data : in   std_logic_vector(7 downto 0);
    input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_data : in   std_logic_vector(7 downto 0);
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(7 downto 0);
    kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_data : in   std_logic_vector(7 downto 0);
    kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_data : in   std_logic_vector(7 downto 0);
    input_pipe4_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe4_pipe_read_data : in   std_logic_vector(7 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(7 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_6623_start: Boolean;
  signal convolve_CP_6623_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_num_out_pipe_2569_inst_ack_1 : boolean;
  signal RPIPE_num_out_pipe_2574_inst_req_1 : boolean;
  signal SUB_u16_u16_2576_inst_ack_0 : boolean;
  signal SUB_u16_u16_2581_inst_req_0 : boolean;
  signal RPIPE_size_pipe_2579_inst_req_1 : boolean;
  signal nacc1_2990_2590_buf_req_0 : boolean;
  signal RPIPE_num_out_pipe_2574_inst_ack_1 : boolean;
  signal SUB_u16_u16_2581_inst_ack_1 : boolean;
  signal SUB_u16_u16_2581_inst_req_1 : boolean;
  signal nacc1_2990_2590_buf_ack_1 : boolean;
  signal RPIPE_num_out_pipe_2574_inst_ack_0 : boolean;
  signal SUB_u16_u16_2576_inst_req_1 : boolean;
  signal SUB_u16_u16_2581_inst_ack_0 : boolean;
  signal SUB_u16_u16_2571_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_2569_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_2574_inst_req_0 : boolean;
  signal SUB_u16_u16_2576_inst_ack_1 : boolean;
  signal SUB_u16_u16_2571_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_2579_inst_ack_1 : boolean;
  signal SUB_u16_u16_2571_inst_req_1 : boolean;
  signal SUB_u16_u16_2571_inst_ack_0 : boolean;
  signal W_num_done_2875_delayed_1_0_2982_inst_ack_1 : boolean;
  signal W_num_done_2881_delayed_1_0_2991_inst_req_0 : boolean;
  signal W_num_done_2881_delayed_1_0_2991_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2927_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2934_inst_req_0 : boolean;
  signal phi_stmt_2585_ack_0 : boolean;
  signal RPIPE_num_out_pipe_2569_inst_ack_0 : boolean;
  signal nacc2_2999_2595_buf_req_0 : boolean;
  signal phi_stmt_2591_req_0 : boolean;
  signal n_row_2981_2600_buf_req_1 : boolean;
  signal phi_stmt_2591_ack_0 : boolean;
  signal nacc2_2999_2595_buf_ack_0 : boolean;
  signal n_row_2981_2600_buf_ack_1 : boolean;
  signal RPIPE_size_pipe_2579_inst_req_0 : boolean;
  signal RPIPE_size_pipe_2579_inst_ack_0 : boolean;
  signal phi_stmt_2601_req_1 : boolean;
  signal W_store_kernel_2824_delayed_1_0_2923_inst_req_1 : boolean;
  signal SUB_u16_u16_2905_inst_req_1 : boolean;
  signal phi_stmt_2585_req_1 : boolean;
  signal do_while_stmt_2583_branch_req_0 : boolean;
  signal W_store_kernel_2824_delayed_1_0_2923_inst_ack_0 : boolean;
  signal phi_stmt_2596_req_1 : boolean;
  signal phi_stmt_2601_ack_0 : boolean;
  signal nacc1_2990_2590_buf_ack_0 : boolean;
  signal nacc2_2999_2595_buf_ack_1 : boolean;
  signal n_row_2981_2600_buf_req_0 : boolean;
  signal W_store_kernel_2824_delayed_1_0_2923_inst_req_0 : boolean;
  signal nacc1_2990_2590_buf_req_1 : boolean;
  signal n_row_2981_2600_buf_ack_0 : boolean;
  signal phi_stmt_2596_ack_0 : boolean;
  signal phi_stmt_2596_req_0 : boolean;
  signal phi_stmt_2591_req_1 : boolean;
  signal phi_stmt_2585_req_0 : boolean;
  signal nacc2_2999_2595_buf_req_1 : boolean;
  signal phi_stmt_2601_req_0 : boolean;
  signal RPIPE_num_out_pipe_2569_inst_req_1 : boolean;
  signal W_store_kernel_2824_delayed_1_0_2923_inst_ack_1 : boolean;
  signal SUB_u16_u16_2576_inst_req_0 : boolean;
  signal W_num_done_2881_delayed_1_0_2991_inst_req_1 : boolean;
  signal W_num_done_2881_delayed_1_0_2991_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2927_inst_ack_0 : boolean;
  signal SUB_u16_u16_2905_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2941_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2941_inst_ack_1 : boolean;
  signal W_store_kernel_2832_delayed_1_0_2937_inst_req_1 : boolean;
  signal W_store_kernel_2832_delayed_1_0_2937_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2934_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2934_inst_ack_1 : boolean;
  signal W_store_kernel_2832_delayed_1_0_2937_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2927_inst_req_1 : boolean;
  signal SUB_u16_u16_2905_inst_req_0 : boolean;
  signal SUB_u16_u16_2905_inst_ack_0 : boolean;
  signal W_num_done_2875_delayed_1_0_2982_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2927_inst_ack_1 : boolean;
  signal W_store_kernel_2828_delayed_1_0_2930_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2941_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2941_inst_ack_0 : boolean;
  signal W_store_kernel_2828_delayed_1_0_2930_inst_ack_0 : boolean;
  signal W_store_kernel_2832_delayed_1_0_2937_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2934_inst_req_1 : boolean;
  signal W_num_done_2875_delayed_1_0_2982_inst_req_0 : boolean;
  signal W_num_done_2875_delayed_1_0_2982_inst_ack_0 : boolean;
  signal W_store_kernel_2828_delayed_1_0_2930_inst_req_1 : boolean;
  signal W_store_kernel_2828_delayed_1_0_2930_inst_ack_1 : boolean;
  signal n_col_2973_2605_buf_req_0 : boolean;
  signal n_col_2973_2605_buf_ack_0 : boolean;
  signal n_col_2973_2605_buf_req_1 : boolean;
  signal n_col_2973_2605_buf_ack_1 : boolean;
  signal phi_stmt_2606_req_1 : boolean;
  signal phi_stmt_2606_req_0 : boolean;
  signal phi_stmt_2606_ack_0 : boolean;
  signal n_num_2962_2611_buf_req_0 : boolean;
  signal n_num_2962_2611_buf_ack_0 : boolean;
  signal n_num_2962_2611_buf_req_1 : boolean;
  signal n_num_2962_2611_buf_ack_1 : boolean;
  signal phi_stmt_2612_req_1 : boolean;
  signal phi_stmt_2612_req_0 : boolean;
  signal phi_stmt_2612_ack_0 : boolean;
  signal n_chl_2951_2616_buf_req_0 : boolean;
  signal n_chl_2951_2616_buf_ack_0 : boolean;
  signal n_chl_2951_2616_buf_req_1 : boolean;
  signal n_chl_2951_2616_buf_ack_1 : boolean;
  signal RPIPE_input_pipe1_2629_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_2629_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_2629_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_2629_inst_ack_1 : boolean;
  signal RPIPE_input_pipe2_2633_inst_req_0 : boolean;
  signal RPIPE_input_pipe2_2633_inst_ack_0 : boolean;
  signal RPIPE_input_pipe2_2633_inst_req_1 : boolean;
  signal RPIPE_input_pipe2_2633_inst_ack_1 : boolean;
  signal RPIPE_input_pipe3_2637_inst_req_0 : boolean;
  signal RPIPE_input_pipe3_2637_inst_ack_0 : boolean;
  signal RPIPE_input_pipe3_2637_inst_req_1 : boolean;
  signal RPIPE_input_pipe3_2637_inst_ack_1 : boolean;
  signal RPIPE_input_pipe4_2641_inst_req_0 : boolean;
  signal RPIPE_input_pipe4_2641_inst_ack_0 : boolean;
  signal RPIPE_input_pipe4_2641_inst_req_1 : boolean;
  signal RPIPE_input_pipe4_2641_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2645_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2645_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2645_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2645_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2649_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2649_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2649_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2649_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2653_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2653_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2653_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2653_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2657_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2657_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2657_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2657_inst_ack_1 : boolean;
  signal W_read_ip_2603_delayed_1_0_2659_inst_req_0 : boolean;
  signal W_read_ip_2603_delayed_1_0_2659_inst_ack_0 : boolean;
  signal W_read_ip_2603_delayed_1_0_2659_inst_req_1 : boolean;
  signal W_read_ip_2603_delayed_1_0_2659_inst_ack_1 : boolean;
  signal W_read_ip_2609_delayed_1_0_2668_inst_req_0 : boolean;
  signal W_read_ip_2609_delayed_1_0_2668_inst_ack_0 : boolean;
  signal W_read_ip_2609_delayed_1_0_2668_inst_req_1 : boolean;
  signal W_read_ip_2609_delayed_1_0_2668_inst_ack_1 : boolean;
  signal W_read_ip_2615_delayed_1_0_2677_inst_req_0 : boolean;
  signal W_read_ip_2615_delayed_1_0_2677_inst_ack_0 : boolean;
  signal W_read_ip_2615_delayed_1_0_2677_inst_req_1 : boolean;
  signal W_read_ip_2615_delayed_1_0_2677_inst_ack_1 : boolean;
  signal W_read_ip_2621_delayed_1_0_2686_inst_req_0 : boolean;
  signal W_read_ip_2621_delayed_1_0_2686_inst_ack_0 : boolean;
  signal W_read_ip_2621_delayed_1_0_2686_inst_req_1 : boolean;
  signal W_read_ip_2621_delayed_1_0_2686_inst_ack_1 : boolean;
  signal W_write_input_2635_delayed_1_0_2704_inst_req_0 : boolean;
  signal W_write_input_2635_delayed_1_0_2704_inst_ack_0 : boolean;
  signal W_write_input_2635_delayed_1_0_2704_inst_req_1 : boolean;
  signal W_write_input_2635_delayed_1_0_2704_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2708_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2708_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2708_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2708_inst_ack_1 : boolean;
  signal W_write_input_2639_delayed_1_0_2711_inst_req_0 : boolean;
  signal W_write_input_2639_delayed_1_0_2711_inst_ack_0 : boolean;
  signal W_write_input_2639_delayed_1_0_2711_inst_req_1 : boolean;
  signal W_write_input_2639_delayed_1_0_2711_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2715_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2715_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2715_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2715_inst_ack_1 : boolean;
  signal W_write_input_2643_delayed_1_0_2718_inst_req_0 : boolean;
  signal W_write_input_2643_delayed_1_0_2718_inst_ack_0 : boolean;
  signal W_write_input_2643_delayed_1_0_2718_inst_req_1 : boolean;
  signal W_write_input_2643_delayed_1_0_2718_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2722_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2722_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2722_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2722_inst_ack_1 : boolean;
  signal W_write_input_2647_delayed_1_0_2725_inst_req_0 : boolean;
  signal W_write_input_2647_delayed_1_0_2725_inst_ack_0 : boolean;
  signal W_write_input_2647_delayed_1_0_2725_inst_req_1 : boolean;
  signal W_write_input_2647_delayed_1_0_2725_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2729_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2729_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2729_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2729_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_2759_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe1_2759_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_2759_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_2759_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe2_2763_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe2_2763_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe2_2763_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe2_2763_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe3_2767_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe3_2767_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe3_2767_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe3_2767_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2771_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2771_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2771_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2771_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2775_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2775_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2775_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2775_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2779_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2779_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2779_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2779_inst_ack_1 : boolean;
  signal W_read_k_2701_delayed_1_0_2781_inst_req_0 : boolean;
  signal W_read_k_2701_delayed_1_0_2781_inst_ack_0 : boolean;
  signal W_read_k_2701_delayed_1_0_2781_inst_req_1 : boolean;
  signal W_read_k_2701_delayed_1_0_2781_inst_ack_1 : boolean;
  signal W_read_k_2707_delayed_1_0_2790_inst_req_0 : boolean;
  signal W_read_k_2707_delayed_1_0_2790_inst_ack_0 : boolean;
  signal W_read_k_2707_delayed_1_0_2790_inst_req_1 : boolean;
  signal W_read_k_2707_delayed_1_0_2790_inst_ack_1 : boolean;
  signal W_read_k_2713_delayed_1_0_2799_inst_req_0 : boolean;
  signal W_read_k_2713_delayed_1_0_2799_inst_ack_0 : boolean;
  signal W_read_k_2713_delayed_1_0_2799_inst_req_1 : boolean;
  signal W_read_k_2713_delayed_1_0_2799_inst_ack_1 : boolean;
  signal W_acc1_2767_delayed_1_0_2856_inst_req_0 : boolean;
  signal W_acc1_2767_delayed_1_0_2856_inst_ack_0 : boolean;
  signal W_acc1_2767_delayed_1_0_2856_inst_req_1 : boolean;
  signal W_acc1_2767_delayed_1_0_2856_inst_ack_1 : boolean;
  signal W_acc2_2776_delayed_1_0_2868_inst_req_0 : boolean;
  signal W_acc2_2776_delayed_1_0_2868_inst_ack_0 : boolean;
  signal W_acc2_2776_delayed_1_0_2868_inst_req_1 : boolean;
  signal W_acc2_2776_delayed_1_0_2868_inst_ack_1 : boolean;
  signal W_num_done_2886_delayed_1_0_3000_inst_req_0 : boolean;
  signal W_num_done_2886_delayed_1_0_3000_inst_ack_0 : boolean;
  signal W_num_done_2886_delayed_1_0_3000_inst_req_1 : boolean;
  signal W_num_done_2886_delayed_1_0_3000_inst_ack_1 : boolean;
  signal CONCAT_u8_u16_3009_inst_req_0 : boolean;
  signal CONCAT_u8_u16_3009_inst_ack_0 : boolean;
  signal CONCAT_u8_u16_3009_inst_req_1 : boolean;
  signal CONCAT_u8_u16_3009_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_3004_inst_req_0 : boolean;
  signal WPIPE_output_pipe_3004_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_3004_inst_req_1 : boolean;
  signal WPIPE_output_pipe_3004_inst_ack_1 : boolean;
  signal do_while_stmt_2583_branch_ack_0 : boolean;
  signal do_while_stmt_2583_branch_ack_1 : boolean;
  signal WPIPE_input_done_pipe_3014_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_3014_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_3014_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_3014_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_6623_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_6623_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_6623_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_6623_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_6623: Block -- control-path 
    signal convolve_CP_6623_elements: BooleanArray(312 downto 0);
    -- 
  begin -- 
    convolve_CP_6623_elements(0) <= convolve_CP_6623_start;
    convolve_CP_6623_symbol <= convolve_CP_6623_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	312 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_2566/branch_block_stmt_2566__entry__
      -- CP-element group 0: 	 branch_block_stmt_2566/merge_stmt_2567__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2566/$entry
      -- CP-element group 0: 	 branch_block_stmt_2566/merge_stmt_2567_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_2566/merge_stmt_2567__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_2566/merge_stmt_2567__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_2566/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2566/branch_block_stmt_2566__exit__
      -- 
    convolve_CP_6623_elements(1) <= false; 
    -- CP-element group 2:  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	309 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	310 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2566/assign_stmt_3016__entry__
      -- CP-element group 2: 	 branch_block_stmt_2566/do_while_stmt_2583__exit__
      -- CP-element group 2: 	 branch_block_stmt_2566/assign_stmt_3016/$entry
      -- CP-element group 2: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_Sample/req
      -- 
    req_7633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(2), ack => WPIPE_input_done_pipe_3014_inst_req_0); -- 
    convolve_CP_6623_elements(2) <= convolve_CP_6623_elements(309);
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	312 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_Update/cr
      -- 
    ra_6655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2569_inst_ack_0, ack => convolve_CP_6623_elements(3)); -- 
    cr_6659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(3), ack => RPIPE_num_out_pipe_2569_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_Sample/$entry
      -- 
    ca_6660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2569_inst_ack_1, ack => convolve_CP_6623_elements(4)); -- 
    rr_6664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(4), ack => SUB_u16_u16_2571_inst_req_0); -- 
    rr_6682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(4), ack => RPIPE_num_out_pipe_2574_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_sample_completed_
      -- 
    ra_6665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2571_inst_ack_0, ack => convolve_CP_6623_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	312 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	15 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_update_completed_
      -- 
    ca_6670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2571_inst_ack_1, ack => convolve_CP_6623_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_update_start_
      -- CP-element group 7: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_Sample/$exit
      -- 
    ra_6683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2574_inst_ack_0, ack => convolve_CP_6623_elements(7)); -- 
    cr_6687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(7), ack => RPIPE_num_out_pipe_2574_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2574_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_Sample/rr
      -- 
    ca_6688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2574_inst_ack_1, ack => convolve_CP_6623_elements(8)); -- 
    rr_6692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(8), ack => SUB_u16_u16_2576_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_Sample/$exit
      -- 
    ra_6693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2576_inst_ack_0, ack => convolve_CP_6623_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	312 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_Update/$exit
      -- 
    ca_6698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2576_inst_ack_1, ack => convolve_CP_6623_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	312 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_update_start_
      -- CP-element group 11: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_Update/$entry
      -- 
    ra_6711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_2579_inst_ack_0, ack => convolve_CP_6623_elements(11)); -- 
    cr_6715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(11), ack => RPIPE_size_pipe_2579_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_Update/$exit
      -- 
    ca_6716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_2579_inst_ack_1, ack => convolve_CP_6623_elements(12)); -- 
    rr_6720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(12), ack => SUB_u16_u16_2581_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_sample_completed_
      -- 
    ra_6721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2581_inst_ack_0, ack => convolve_CP_6623_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	312 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_Update/$exit
      -- 
    ca_6726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2581_inst_ack_1, ack => convolve_CP_6623_elements(14)); -- 
    -- CP-element group 15:  join  transition  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	6 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582__exit__
      -- CP-element group 15: 	 branch_block_stmt_2566/do_while_stmt_2583__entry__
      -- CP-element group 15: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/$exit
      -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(14) & convolve_CP_6623_elements(10) & convolve_CP_6623_elements(6);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583__entry__
      -- CP-element group 16: 	 branch_block_stmt_2566/do_while_stmt_2583/$entry
      -- 
    convolve_CP_6623_elements(16) <= convolve_CP_6623_elements(15);
    -- CP-element group 17:  merge  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	309 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583__exit__
      -- 
    -- Element group convolve_CP_6623_elements(17) is bound as output of CP function.
    -- CP-element group 18:  merge  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2566/do_while_stmt_2583/loop_back
      -- 
    -- Element group convolve_CP_6623_elements(18) is bound as output of CP function.
    -- CP-element group 19:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	307 
    -- CP-element group 19: 	308 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2566/do_while_stmt_2583/condition_done
      -- CP-element group 19: 	 branch_block_stmt_2566/do_while_stmt_2583/loop_exit/$entry
      -- CP-element group 19: 	 branch_block_stmt_2566/do_while_stmt_2583/loop_taken/$entry
      -- 
    convolve_CP_6623_elements(19) <= convolve_CP_6623_elements(24);
    -- CP-element group 20:  branch  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	306 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2566/do_while_stmt_2583/loop_body_done
      -- 
    convolve_CP_6623_elements(20) <= convolve_CP_6623_elements(306);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	33 
    -- CP-element group 21: 	52 
    -- CP-element group 21: 	71 
    -- CP-element group 21: 	90 
    -- CP-element group 21: 	128 
    -- CP-element group 21: 	109 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_6623_elements(21) <= convolve_CP_6623_elements(18);
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	35 
    -- CP-element group 22: 	54 
    -- CP-element group 22: 	73 
    -- CP-element group 22: 	92 
    -- CP-element group 22: 	130 
    -- CP-element group 22: 	111 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_6623_elements(22) <= convolve_CP_6623_elements(16);
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	225 
    -- CP-element group 23: 	229 
    -- CP-element group 23: 	233 
    -- CP-element group 23: 	237 
    -- CP-element group 23: 	217 
    -- CP-element group 23: 	221 
    -- CP-element group 23: 	161 
    -- CP-element group 23: 	165 
    -- CP-element group 23: 	29 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	46 
    -- CP-element group 23: 	47 
    -- CP-element group 23: 	65 
    -- CP-element group 23: 	66 
    -- CP-element group 23: 	84 
    -- CP-element group 23: 	85 
    -- CP-element group 23: 	169 
    -- CP-element group 23: 	157 
    -- CP-element group 23: 	122 
    -- CP-element group 23: 	123 
    -- CP-element group 23: 	103 
    -- CP-element group 23: 	104 
    -- CP-element group 23: 	261 
    -- CP-element group 23: 	141 
    -- CP-element group 23: 	145 
    -- CP-element group 23: 	149 
    -- CP-element group 23: 	153 
    -- CP-element group 23: 	305 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/$entry
      -- CP-element group 23: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_6623_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	70 
    -- CP-element group 24: 	89 
    -- CP-element group 24: 	127 
    -- CP-element group 24: 	108 
    -- CP-element group 24: 	264 
    -- CP-element group 24: 	305 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	19 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/condition_evaluated
      -- 
    condition_evaluated_6741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_6741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(24), ack => do_while_stmt_2583_branch_req_0); -- 
    convolve_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(28) & convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(127) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(264) & convolve_CP_6623_elements(305);
      gj_convolve_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	29 
    -- CP-element group 25: 	46 
    -- CP-element group 25: 	65 
    -- CP-element group 25: 	84 
    -- CP-element group 25: 	122 
    -- CP-element group 25: 	103 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	28 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	48 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	86 
    -- CP-element group 25: 	124 
    -- CP-element group 25: 	105 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/aggregated_phi_sample_req
      -- 
    convolve_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(29) & convolve_CP_6623_elements(46) & convolve_CP_6623_elements(65) & convolve_CP_6623_elements(84) & convolve_CP_6623_elements(122) & convolve_CP_6623_elements(103) & convolve_CP_6623_elements(28);
      gj_convolve_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: 	49 
    -- CP-element group 26: 	68 
    -- CP-element group 26: 	87 
    -- CP-element group 26: 	125 
    -- CP-element group 26: 	106 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	226 
    -- CP-element group 26: 	230 
    -- CP-element group 26: 	234 
    -- CP-element group 26: 	238 
    -- CP-element group 26: 	218 
    -- CP-element group 26: 	222 
    -- CP-element group 26: 	162 
    -- CP-element group 26: 	166 
    -- CP-element group 26: 	170 
    -- CP-element group 26: 	154 
    -- CP-element group 26: 	158 
    -- CP-element group 26: 	182 
    -- CP-element group 26: 	186 
    -- CP-element group 26: 	254 
    -- CP-element group 26: 	258 
    -- CP-element group 26: 	142 
    -- CP-element group 26: 	146 
    -- CP-element group 26: 	150 
    -- CP-element group 26: 	242 
    -- CP-element group 26: 	246 
    -- CP-element group 26: 	250 
    -- CP-element group 26: 	174 
    -- CP-element group 26: 	178 
    -- CP-element group 26: 	287 
    -- CP-element group 26: 	291 
    -- CP-element group 26: 	306 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26: 	46 
    -- CP-element group 26: 	65 
    -- CP-element group 26: 	84 
    -- CP-element group 26: 	122 
    -- CP-element group 26: 	103 
    -- CP-element group 26:  members (7) 
      -- CP-element group 26: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/aggregated_phi_sample_ack
      -- CP-element group 26: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_sample_completed_
      -- 
    convolve_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(31) & convolve_CP_6623_elements(49) & convolve_CP_6623_elements(68) & convolve_CP_6623_elements(87) & convolve_CP_6623_elements(125) & convolve_CP_6623_elements(106);
      gj_convolve_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	47 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	85 
    -- CP-element group 27: 	123 
    -- CP-element group 27: 	104 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	50 
    -- CP-element group 27: 	69 
    -- CP-element group 27: 	88 
    -- CP-element group 27: 	126 
    -- CP-element group 27: 	107 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/aggregated_phi_update_req
      -- 
    convolve_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(30) & convolve_CP_6623_elements(47) & convolve_CP_6623_elements(66) & convolve_CP_6623_elements(85) & convolve_CP_6623_elements(123) & convolve_CP_6623_elements(104);
      gj_convolve_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	32 
    -- CP-element group 28: 	51 
    -- CP-element group 28: 	70 
    -- CP-element group 28: 	89 
    -- CP-element group 28: 	127 
    -- CP-element group 28: 	108 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	25 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(32) & convolve_CP_6623_elements(51) & convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(127) & convolve_CP_6623_elements(108);
      gj_convolve_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	224 
    -- CP-element group 29: 	228 
    -- CP-element group 29: 	232 
    -- CP-element group 29: 	236 
    -- CP-element group 29: 	220 
    -- CP-element group 29: 	160 
    -- CP-element group 29: 	164 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	168 
    -- CP-element group 29: 	180 
    -- CP-element group 29: 	184 
    -- CP-element group 29: 	256 
    -- CP-element group 29: 	144 
    -- CP-element group 29: 	148 
    -- CP-element group 29: 	152 
    -- CP-element group 29: 	240 
    -- CP-element group 29: 	244 
    -- CP-element group 29: 	248 
    -- CP-element group 29: 	252 
    -- CP-element group 29: 	176 
    -- CP-element group 29: 	289 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_sample_start_
      -- 
    convolve_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(224) & convolve_CP_6623_elements(228) & convolve_CP_6623_elements(232) & convolve_CP_6623_elements(236) & convolve_CP_6623_elements(220) & convolve_CP_6623_elements(160) & convolve_CP_6623_elements(164) & convolve_CP_6623_elements(26) & convolve_CP_6623_elements(168) & convolve_CP_6623_elements(180) & convolve_CP_6623_elements(184) & convolve_CP_6623_elements(256) & convolve_CP_6623_elements(144) & convolve_CP_6623_elements(148) & convolve_CP_6623_elements(152) & convolve_CP_6623_elements(240) & convolve_CP_6623_elements(244) & convolve_CP_6623_elements(248) & convolve_CP_6623_elements(252) & convolve_CP_6623_elements(176) & convolve_CP_6623_elements(289);
      gj_convolve_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	23 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	255 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	27 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_update_start_
      -- 
    convolve_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(32) & convolve_CP_6623_elements(255);
      gj_convolve_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	26 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_sample_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(31) is bound as output of CP function.
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	28 
    -- CP-element group 32: 	253 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_update_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(32) is bound as output of CP function.
    -- CP-element group 33:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	21 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_loopback_trigger
      -- 
    convolve_CP_6623_elements(33) <= convolve_CP_6623_elements(21);
    -- CP-element group 34:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_loopback_sample_req
      -- CP-element group 34: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_loopback_sample_req_ps
      -- 
    phi_stmt_2585_loopback_sample_req_6756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2585_loopback_sample_req_6756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(34), ack => phi_stmt_2585_req_1); -- 
    -- Element group convolve_CP_6623_elements(34) is bound as output of CP function.
    -- CP-element group 35:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	22 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_entry_trigger
      -- 
    convolve_CP_6623_elements(35) <= convolve_CP_6623_elements(22);
    -- CP-element group 36:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_entry_sample_req
      -- CP-element group 36: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_entry_sample_req_ps
      -- 
    phi_stmt_2585_entry_sample_req_6759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2585_entry_sample_req_6759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(36), ack => phi_stmt_2585_req_0); -- 
    -- Element group convolve_CP_6623_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_phi_mux_ack_ps
      -- CP-element group 37: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2585_phi_mux_ack
      -- 
    phi_stmt_2585_phi_mux_ack_6762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2585_ack_0, ack => convolve_CP_6623_elements(37)); -- 
    -- CP-element group 38:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2589_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2589_sample_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2589_sample_start__ps
      -- CP-element group 38: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2589_sample_completed_
      -- 
    -- Element group convolve_CP_6623_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2589_update_start__ps
      -- CP-element group 39: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2589_update_start_
      -- 
    -- Element group convolve_CP_6623_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2589_update_completed__ps
      -- 
    convolve_CP_6623_elements(40) <= convolve_CP_6623_elements(41);
    -- CP-element group 41:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	40 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2589_update_completed_
      -- 
    -- Element group convolve_CP_6623_elements(41) is a control-delay.
    cp_element_41_delay: control_delay_element  generic map(name => " 41_delay", delay_value => 1)  port map(req => convolve_CP_6623_elements(39), ack => convolve_CP_6623_elements(41), clk => clk, reset =>reset);
    -- CP-element group 42:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_Sample/req
      -- CP-element group 42: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_sample_start__ps
      -- CP-element group 42: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_sample_start_
      -- 
    req_6783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(42), ack => nacc1_2990_2590_buf_req_0); -- 
    -- Element group convolve_CP_6623_elements(42) is bound as output of CP function.
    -- CP-element group 43:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_update_start_
      -- CP-element group 43: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_update_start__ps
      -- CP-element group 43: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_Update/req
      -- 
    req_6788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(43), ack => nacc1_2990_2590_buf_req_1); -- 
    -- Element group convolve_CP_6623_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_sample_completed__ps
      -- CP-element group 44: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_Sample/ack
      -- 
    ack_6784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc1_2990_2590_buf_ack_0, ack => convolve_CP_6623_elements(44)); -- 
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_Update/ack
      -- CP-element group 45: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_update_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc1_2590_Update/$exit
      -- 
    ack_6789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc1_2990_2590_buf_ack_1, ack => convolve_CP_6623_elements(45)); -- 
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	224 
    -- CP-element group 46: 	228 
    -- CP-element group 46: 	232 
    -- CP-element group 46: 	236 
    -- CP-element group 46: 	220 
    -- CP-element group 46: 	164 
    -- CP-element group 46: 	26 
    -- CP-element group 46: 	168 
    -- CP-element group 46: 	172 
    -- CP-element group 46: 	156 
    -- CP-element group 46: 	180 
    -- CP-element group 46: 	184 
    -- CP-element group 46: 	188 
    -- CP-element group 46: 	260 
    -- CP-element group 46: 	148 
    -- CP-element group 46: 	152 
    -- CP-element group 46: 	240 
    -- CP-element group 46: 	244 
    -- CP-element group 46: 	248 
    -- CP-element group 46: 	252 
    -- CP-element group 46: 	293 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	25 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_sample_start_
      -- 
    convolve_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(224) & convolve_CP_6623_elements(228) & convolve_CP_6623_elements(232) & convolve_CP_6623_elements(236) & convolve_CP_6623_elements(220) & convolve_CP_6623_elements(164) & convolve_CP_6623_elements(26) & convolve_CP_6623_elements(168) & convolve_CP_6623_elements(172) & convolve_CP_6623_elements(156) & convolve_CP_6623_elements(180) & convolve_CP_6623_elements(184) & convolve_CP_6623_elements(188) & convolve_CP_6623_elements(260) & convolve_CP_6623_elements(148) & convolve_CP_6623_elements(152) & convolve_CP_6623_elements(240) & convolve_CP_6623_elements(244) & convolve_CP_6623_elements(248) & convolve_CP_6623_elements(252) & convolve_CP_6623_elements(293);
      gj_convolve_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	23 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	51 
    -- CP-element group 47: 	259 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	27 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_update_start_
      -- 
    convolve_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(51) & convolve_CP_6623_elements(259);
      gj_convolve_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	25 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_sample_start__ps
      -- 
    convolve_CP_6623_elements(48) <= convolve_CP_6623_elements(25);
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	26 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_sample_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(49) is bound as output of CP function.
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	27 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_update_start__ps
      -- 
    convolve_CP_6623_elements(50) <= convolve_CP_6623_elements(27);
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	28 
    -- CP-element group 51: 	257 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	47 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_update_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	21 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_loopback_trigger
      -- 
    convolve_CP_6623_elements(52) <= convolve_CP_6623_elements(21);
    -- CP-element group 53:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_loopback_sample_req_ps
      -- CP-element group 53: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_loopback_sample_req
      -- 
    phi_stmt_2591_loopback_sample_req_6800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2591_loopback_sample_req_6800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(53), ack => phi_stmt_2591_req_1); -- 
    -- Element group convolve_CP_6623_elements(53) is bound as output of CP function.
    -- CP-element group 54:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	22 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_entry_trigger
      -- 
    convolve_CP_6623_elements(54) <= convolve_CP_6623_elements(22);
    -- CP-element group 55:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_entry_sample_req
      -- CP-element group 55: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_entry_sample_req_ps
      -- 
    phi_stmt_2591_entry_sample_req_6803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2591_entry_sample_req_6803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(55), ack => phi_stmt_2591_req_0); -- 
    -- Element group convolve_CP_6623_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_phi_mux_ack_ps
      -- CP-element group 56: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2591_phi_mux_ack
      -- 
    phi_stmt_2591_phi_mux_ack_6806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2591_ack_0, ack => convolve_CP_6623_elements(56)); -- 
    -- CP-element group 57:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2594_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2594_sample_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2594_sample_start__ps
      -- CP-element group 57: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2594_sample_completed_
      -- 
    -- Element group convolve_CP_6623_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2594_update_start_
      -- CP-element group 58: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2594_update_start__ps
      -- 
    -- Element group convolve_CP_6623_elements(58) is bound as output of CP function.
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2594_update_completed__ps
      -- 
    convolve_CP_6623_elements(59) <= convolve_CP_6623_elements(60);
    -- CP-element group 60:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	59 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2594_update_completed_
      -- 
    -- Element group convolve_CP_6623_elements(60) is a control-delay.
    cp_element_60_delay: control_delay_element  generic map(name => " 60_delay", delay_value => 1)  port map(req => convolve_CP_6623_elements(58), ack => convolve_CP_6623_elements(60), clk => clk, reset =>reset);
    -- CP-element group 61:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_sample_start__ps
      -- CP-element group 61: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_Sample/req
      -- CP-element group 61: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_sample_start_
      -- 
    req_6827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(61), ack => nacc2_2999_2595_buf_req_0); -- 
    -- Element group convolve_CP_6623_elements(61) is bound as output of CP function.
    -- CP-element group 62:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_update_start__ps
      -- CP-element group 62: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_Update/req
      -- CP-element group 62: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_update_start_
      -- 
    req_6832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(62), ack => nacc2_2999_2595_buf_req_1); -- 
    -- Element group convolve_CP_6623_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_sample_completed__ps
      -- CP-element group 63: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_sample_completed_
      -- 
    ack_6828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc2_2999_2595_buf_ack_0, ack => convolve_CP_6623_elements(63)); -- 
    -- CP-element group 64:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_update_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_nacc2_2595_Update/$exit
      -- 
    ack_6833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc2_2999_2595_buf_ack_1, ack => convolve_CP_6623_elements(64)); -- 
    -- CP-element group 65:  join  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	23 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	26 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	25 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_sample_start_
      -- 
    convolve_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(26);
      gj_convolve_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  join  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	23 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	226 
    -- CP-element group 66: 	230 
    -- CP-element group 66: 	234 
    -- CP-element group 66: 	238 
    -- CP-element group 66: 	218 
    -- CP-element group 66: 	222 
    -- CP-element group 66: 	70 
    -- CP-element group 66: 	243 
    -- CP-element group 66: 	247 
    -- CP-element group 66: 	251 
    -- CP-element group 66: 	267 
    -- CP-element group 66: 	274 
    -- CP-element group 66: 	281 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	27 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_update_start_
      -- 
    convolve_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(226) & convolve_CP_6623_elements(230) & convolve_CP_6623_elements(234) & convolve_CP_6623_elements(238) & convolve_CP_6623_elements(218) & convolve_CP_6623_elements(222) & convolve_CP_6623_elements(70) & convolve_CP_6623_elements(243) & convolve_CP_6623_elements(247) & convolve_CP_6623_elements(251) & convolve_CP_6623_elements(267) & convolve_CP_6623_elements(274) & convolve_CP_6623_elements(281);
      gj_convolve_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_sample_start__ps
      -- 
    convolve_CP_6623_elements(67) <= convolve_CP_6623_elements(25);
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	26 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_sample_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(68) is bound as output of CP function.
    -- CP-element group 69:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	27 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_update_start__ps
      -- 
    convolve_CP_6623_elements(69) <= convolve_CP_6623_elements(27);
    -- CP-element group 70:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	226 
    -- CP-element group 70: 	230 
    -- CP-element group 70: 	234 
    -- CP-element group 70: 	238 
    -- CP-element group 70: 	218 
    -- CP-element group 70: 	222 
    -- CP-element group 70: 	24 
    -- CP-element group 70: 	28 
    -- CP-element group 70: 	265 
    -- CP-element group 70: 	241 
    -- CP-element group 70: 	245 
    -- CP-element group 70: 	249 
    -- CP-element group 70: 	272 
    -- CP-element group 70: 	279 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	66 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_update_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(70) is bound as output of CP function.
    -- CP-element group 71:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	21 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_loopback_trigger
      -- 
    convolve_CP_6623_elements(71) <= convolve_CP_6623_elements(21);
    -- CP-element group 72:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_loopback_sample_req
      -- CP-element group 72: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_loopback_sample_req_ps
      -- 
    phi_stmt_2596_loopback_sample_req_6844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2596_loopback_sample_req_6844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(72), ack => phi_stmt_2596_req_1); -- 
    -- Element group convolve_CP_6623_elements(72) is bound as output of CP function.
    -- CP-element group 73:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	22 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_entry_trigger
      -- 
    convolve_CP_6623_elements(73) <= convolve_CP_6623_elements(22);
    -- CP-element group 74:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_entry_sample_req
      -- CP-element group 74: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_entry_sample_req_ps
      -- 
    phi_stmt_2596_entry_sample_req_6847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2596_entry_sample_req_6847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(74), ack => phi_stmt_2596_req_0); -- 
    -- Element group convolve_CP_6623_elements(74) is bound as output of CP function.
    -- CP-element group 75:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_phi_mux_ack
      -- CP-element group 75: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2596_phi_mux_ack_ps
      -- 
    phi_stmt_2596_phi_mux_ack_6850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2596_ack_0, ack => convolve_CP_6623_elements(75)); -- 
    -- CP-element group 76:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2599_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2599_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2599_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2599_sample_start__ps
      -- 
    -- Element group convolve_CP_6623_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2599_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2599_update_start__ps
      -- 
    -- Element group convolve_CP_6623_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2599_update_completed__ps
      -- 
    convolve_CP_6623_elements(78) <= convolve_CP_6623_elements(79);
    -- CP-element group 79:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	78 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2599_update_completed_
      -- 
    -- Element group convolve_CP_6623_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convolve_CP_6623_elements(77), ack => convolve_CP_6623_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_Sample/req
      -- CP-element group 80: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_sample_start__ps
      -- 
    req_6871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(80), ack => n_row_2981_2600_buf_req_0); -- 
    -- Element group convolve_CP_6623_elements(80) is bound as output of CP function.
    -- CP-element group 81:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_update_start_
      -- CP-element group 81: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_Update/req
      -- CP-element group 81: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_update_start__ps
      -- 
    req_6876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(81), ack => n_row_2981_2600_buf_req_1); -- 
    -- Element group convolve_CP_6623_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_sample_completed__ps
      -- CP-element group 82: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_Sample/ack
      -- 
    ack_6872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_2981_2600_buf_ack_0, ack => convolve_CP_6623_elements(82)); -- 
    -- CP-element group 83:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_Update/ack
      -- CP-element group 83: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_row_2600_update_completed__ps
      -- 
    ack_6877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_2981_2600_buf_ack_1, ack => convolve_CP_6623_elements(83)); -- 
    -- CP-element group 84:  join  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	23 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	26 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	25 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_sample_start_
      -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(26);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	23 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	226 
    -- CP-element group 85: 	230 
    -- CP-element group 85: 	234 
    -- CP-element group 85: 	238 
    -- CP-element group 85: 	212 
    -- CP-element group 85: 	198 
    -- CP-element group 85: 	218 
    -- CP-element group 85: 	222 
    -- CP-element group 85: 	162 
    -- CP-element group 85: 	166 
    -- CP-element group 85: 	89 
    -- CP-element group 85: 	170 
    -- CP-element group 85: 	154 
    -- CP-element group 85: 	158 
    -- CP-element group 85: 	183 
    -- CP-element group 85: 	187 
    -- CP-element group 85: 	191 
    -- CP-element group 85: 	142 
    -- CP-element group 85: 	146 
    -- CP-element group 85: 	150 
    -- CP-element group 85: 	205 
    -- CP-element group 85: 	243 
    -- CP-element group 85: 	247 
    -- CP-element group 85: 	251 
    -- CP-element group 85: 	175 
    -- CP-element group 85: 	179 
    -- CP-element group 85: 	267 
    -- CP-element group 85: 	274 
    -- CP-element group 85: 	281 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	27 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_update_start_
      -- 
    convolve_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 29) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1);
      constant place_markings: IntegerArray(0 to 29)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1);
      constant place_delays: IntegerArray(0 to 29) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 30); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(226) & convolve_CP_6623_elements(230) & convolve_CP_6623_elements(234) & convolve_CP_6623_elements(238) & convolve_CP_6623_elements(212) & convolve_CP_6623_elements(198) & convolve_CP_6623_elements(218) & convolve_CP_6623_elements(222) & convolve_CP_6623_elements(162) & convolve_CP_6623_elements(166) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(170) & convolve_CP_6623_elements(154) & convolve_CP_6623_elements(158) & convolve_CP_6623_elements(183) & convolve_CP_6623_elements(187) & convolve_CP_6623_elements(191) & convolve_CP_6623_elements(142) & convolve_CP_6623_elements(146) & convolve_CP_6623_elements(150) & convolve_CP_6623_elements(205) & convolve_CP_6623_elements(243) & convolve_CP_6623_elements(247) & convolve_CP_6623_elements(251) & convolve_CP_6623_elements(175) & convolve_CP_6623_elements(179) & convolve_CP_6623_elements(267) & convolve_CP_6623_elements(274) & convolve_CP_6623_elements(281);
      gj_convolve_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 30, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	25 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_sample_start__ps
      -- 
    convolve_CP_6623_elements(86) <= convolve_CP_6623_elements(25);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	26 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_sample_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(87) is bound as output of CP function.
    -- CP-element group 88:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	27 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_update_start__ps
      -- 
    convolve_CP_6623_elements(88) <= convolve_CP_6623_elements(27);
    -- CP-element group 89:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	226 
    -- CP-element group 89: 	230 
    -- CP-element group 89: 	234 
    -- CP-element group 89: 	238 
    -- CP-element group 89: 	210 
    -- CP-element group 89: 	196 
    -- CP-element group 89: 	218 
    -- CP-element group 89: 	222 
    -- CP-element group 89: 	162 
    -- CP-element group 89: 	166 
    -- CP-element group 89: 	24 
    -- CP-element group 89: 	28 
    -- CP-element group 89: 	203 
    -- CP-element group 89: 	170 
    -- CP-element group 89: 	173 
    -- CP-element group 89: 	154 
    -- CP-element group 89: 	158 
    -- CP-element group 89: 	181 
    -- CP-element group 89: 	185 
    -- CP-element group 89: 	189 
    -- CP-element group 89: 	265 
    -- CP-element group 89: 	142 
    -- CP-element group 89: 	146 
    -- CP-element group 89: 	150 
    -- CP-element group 89: 	241 
    -- CP-element group 89: 	245 
    -- CP-element group 89: 	249 
    -- CP-element group 89: 	177 
    -- CP-element group 89: 	272 
    -- CP-element group 89: 	279 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	85 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_update_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_update_completed_
      -- 
    -- Element group convolve_CP_6623_elements(89) is bound as output of CP function.
    -- CP-element group 90:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	21 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_loopback_trigger
      -- 
    convolve_CP_6623_elements(90) <= convolve_CP_6623_elements(21);
    -- CP-element group 91:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_loopback_sample_req
      -- CP-element group 91: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_loopback_sample_req_ps
      -- 
    phi_stmt_2601_loopback_sample_req_6888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2601_loopback_sample_req_6888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(91), ack => phi_stmt_2601_req_1); -- 
    -- Element group convolve_CP_6623_elements(91) is bound as output of CP function.
    -- CP-element group 92:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	22 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_entry_trigger
      -- 
    convolve_CP_6623_elements(92) <= convolve_CP_6623_elements(22);
    -- CP-element group 93:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_entry_sample_req_ps
      -- CP-element group 93: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_entry_sample_req
      -- 
    phi_stmt_2601_entry_sample_req_6891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2601_entry_sample_req_6891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(93), ack => phi_stmt_2601_req_0); -- 
    -- Element group convolve_CP_6623_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_phi_mux_ack
      -- CP-element group 94: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2601_phi_mux_ack_ps
      -- 
    phi_stmt_2601_phi_mux_ack_6894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2601_ack_0, ack => convolve_CP_6623_elements(94)); -- 
    -- CP-element group 95:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2604_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2604_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2604_sample_start__ps
      -- CP-element group 95: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2604_sample_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(95) is bound as output of CP function.
    -- CP-element group 96:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2604_update_start__ps
      -- CP-element group 96: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2604_update_start_
      -- 
    -- Element group convolve_CP_6623_elements(96) is bound as output of CP function.
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2604_update_completed__ps
      -- 
    convolve_CP_6623_elements(97) <= convolve_CP_6623_elements(98);
    -- CP-element group 98:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	97 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2604_update_completed_
      -- 
    -- Element group convolve_CP_6623_elements(98) is a control-delay.
    cp_element_98_delay: control_delay_element  generic map(name => " 98_delay", delay_value => 1)  port map(req => convolve_CP_6623_elements(96), ack => convolve_CP_6623_elements(98), clk => clk, reset =>reset);
    -- CP-element group 99:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (4) 
      -- CP-element group 99: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_sample_start__ps
      -- CP-element group 99: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_Sample/req
      -- 
    req_6915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(99), ack => n_col_2973_2605_buf_req_0); -- 
    -- Element group convolve_CP_6623_elements(99) is bound as output of CP function.
    -- CP-element group 100:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_update_start__ps
      -- CP-element group 100: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_Update/req
      -- 
    req_6920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(100), ack => n_col_2973_2605_buf_req_1); -- 
    -- Element group convolve_CP_6623_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_sample_completed__ps
      -- CP-element group 101: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_Sample/ack
      -- 
    ack_6916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_2973_2605_buf_ack_0, ack => convolve_CP_6623_elements(101)); -- 
    -- CP-element group 102:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_update_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_col_2605_Update/ack
      -- 
    ack_6921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_2973_2605_buf_ack_1, ack => convolve_CP_6623_elements(102)); -- 
    -- CP-element group 103:  join  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	23 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	26 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	25 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_sample_start_
      -- 
    convolve_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(26);
      gj_convolve_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	23 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	212 
    -- CP-element group 104: 	198 
    -- CP-element group 104: 	162 
    -- CP-element group 104: 	166 
    -- CP-element group 104: 	170 
    -- CP-element group 104: 	154 
    -- CP-element group 104: 	158 
    -- CP-element group 104: 	183 
    -- CP-element group 104: 	187 
    -- CP-element group 104: 	191 
    -- CP-element group 104: 	108 
    -- CP-element group 104: 	142 
    -- CP-element group 104: 	146 
    -- CP-element group 104: 	150 
    -- CP-element group 104: 	205 
    -- CP-element group 104: 	175 
    -- CP-element group 104: 	179 
    -- CP-element group 104: 	288 
    -- CP-element group 104: 	292 
    -- CP-element group 104: 	296 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	27 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_update_start_
      -- 
    convolve_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(212) & convolve_CP_6623_elements(198) & convolve_CP_6623_elements(162) & convolve_CP_6623_elements(166) & convolve_CP_6623_elements(170) & convolve_CP_6623_elements(154) & convolve_CP_6623_elements(158) & convolve_CP_6623_elements(183) & convolve_CP_6623_elements(187) & convolve_CP_6623_elements(191) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(142) & convolve_CP_6623_elements(146) & convolve_CP_6623_elements(150) & convolve_CP_6623_elements(205) & convolve_CP_6623_elements(175) & convolve_CP_6623_elements(179) & convolve_CP_6623_elements(288) & convolve_CP_6623_elements(292) & convolve_CP_6623_elements(296);
      gj_convolve_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	25 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_sample_start__ps
      -- 
    convolve_CP_6623_elements(105) <= convolve_CP_6623_elements(25);
    -- CP-element group 106:  join  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	26 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_sample_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(106) is bound as output of CP function.
    -- CP-element group 107:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	27 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_update_start__ps
      -- 
    convolve_CP_6623_elements(107) <= convolve_CP_6623_elements(27);
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	210 
    -- CP-element group 108: 	196 
    -- CP-element group 108: 	162 
    -- CP-element group 108: 	166 
    -- CP-element group 108: 	24 
    -- CP-element group 108: 	28 
    -- CP-element group 108: 	203 
    -- CP-element group 108: 	170 
    -- CP-element group 108: 	173 
    -- CP-element group 108: 	154 
    -- CP-element group 108: 	158 
    -- CP-element group 108: 	181 
    -- CP-element group 108: 	185 
    -- CP-element group 108: 	189 
    -- CP-element group 108: 	142 
    -- CP-element group 108: 	146 
    -- CP-element group 108: 	150 
    -- CP-element group 108: 	177 
    -- CP-element group 108: 	286 
    -- CP-element group 108: 	290 
    -- CP-element group 108: 	294 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	104 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_update_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(108) is bound as output of CP function.
    -- CP-element group 109:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	21 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_loopback_trigger
      -- 
    convolve_CP_6623_elements(109) <= convolve_CP_6623_elements(21);
    -- CP-element group 110:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_loopback_sample_req
      -- CP-element group 110: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_loopback_sample_req_ps
      -- 
    phi_stmt_2606_loopback_sample_req_6932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2606_loopback_sample_req_6932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(110), ack => phi_stmt_2606_req_1); -- 
    -- Element group convolve_CP_6623_elements(110) is bound as output of CP function.
    -- CP-element group 111:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	22 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_entry_trigger
      -- 
    convolve_CP_6623_elements(111) <= convolve_CP_6623_elements(22);
    -- CP-element group 112:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_entry_sample_req
      -- CP-element group 112: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_entry_sample_req_ps
      -- 
    phi_stmt_2606_entry_sample_req_6935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2606_entry_sample_req_6935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(112), ack => phi_stmt_2606_req_0); -- 
    -- Element group convolve_CP_6623_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_phi_mux_ack
      -- CP-element group 113: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2606_phi_mux_ack_ps
      -- 
    phi_stmt_2606_phi_mux_ack_6938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2606_ack_0, ack => convolve_CP_6623_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2610_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2610_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2610_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2610_sample_completed_
      -- 
    -- Element group convolve_CP_6623_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2610_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2610_update_start_
      -- 
    -- Element group convolve_CP_6623_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2610_update_completed__ps
      -- 
    convolve_CP_6623_elements(116) <= convolve_CP_6623_elements(117);
    -- CP-element group 117:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2610_update_completed_
      -- 
    -- Element group convolve_CP_6623_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => convolve_CP_6623_elements(115), ack => convolve_CP_6623_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_sample_start__ps
      -- CP-element group 118: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_Sample/req
      -- 
    req_6959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(118), ack => n_num_2962_2611_buf_req_0); -- 
    -- Element group convolve_CP_6623_elements(118) is bound as output of CP function.
    -- CP-element group 119:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_update_start__ps
      -- CP-element group 119: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_update_start_
      -- CP-element group 119: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_Update/req
      -- 
    req_6964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(119), ack => n_num_2962_2611_buf_req_1); -- 
    -- Element group convolve_CP_6623_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (4) 
      -- CP-element group 120: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_sample_completed__ps
      -- CP-element group 120: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_Sample/ack
      -- 
    ack_6960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_2962_2611_buf_ack_0, ack => convolve_CP_6623_elements(120)); -- 
    -- CP-element group 121:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_update_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_num_2611_Update/ack
      -- 
    ack_6965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_2962_2611_buf_ack_1, ack => convolve_CP_6623_elements(121)); -- 
    -- CP-element group 122:  join  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	23 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	26 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	25 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_sample_start_
      -- 
    convolve_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(26);
      gj_convolve_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	23 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	127 
    -- CP-element group 123: 	288 
    -- CP-element group 123: 	292 
    -- CP-element group 123: 	296 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	27 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_update_start_
      -- 
    convolve_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(127) & convolve_CP_6623_elements(288) & convolve_CP_6623_elements(292) & convolve_CP_6623_elements(296);
      gj_convolve_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	25 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_sample_start__ps
      -- 
    convolve_CP_6623_elements(124) <= convolve_CP_6623_elements(25);
    -- CP-element group 125:  join  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	26 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_sample_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	27 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_update_start__ps
      -- 
    convolve_CP_6623_elements(126) <= convolve_CP_6623_elements(27);
    -- CP-element group 127:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	24 
    -- CP-element group 127: 	28 
    -- CP-element group 127: 	286 
    -- CP-element group 127: 	290 
    -- CP-element group 127: 	294 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	123 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_update_completed__ps
      -- 
    -- Element group convolve_CP_6623_elements(127) is bound as output of CP function.
    -- CP-element group 128:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	21 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_loopback_trigger
      -- 
    convolve_CP_6623_elements(128) <= convolve_CP_6623_elements(21);
    -- CP-element group 129:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_loopback_sample_req
      -- CP-element group 129: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_loopback_sample_req_ps
      -- 
    phi_stmt_2612_loopback_sample_req_6976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2612_loopback_sample_req_6976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(129), ack => phi_stmt_2612_req_1); -- 
    -- Element group convolve_CP_6623_elements(129) is bound as output of CP function.
    -- CP-element group 130:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	22 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_entry_trigger
      -- 
    convolve_CP_6623_elements(130) <= convolve_CP_6623_elements(22);
    -- CP-element group 131:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_entry_sample_req
      -- CP-element group 131: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_entry_sample_req_ps
      -- 
    phi_stmt_2612_entry_sample_req_6979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2612_entry_sample_req_6979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(131), ack => phi_stmt_2612_req_0); -- 
    -- Element group convolve_CP_6623_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_phi_mux_ack
      -- CP-element group 132: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/phi_stmt_2612_phi_mux_ack_ps
      -- 
    phi_stmt_2612_phi_mux_ack_6982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2612_ack_0, ack => convolve_CP_6623_elements(132)); -- 
    -- CP-element group 133:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2615_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2615_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2615_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2615_sample_completed_
      -- 
    -- Element group convolve_CP_6623_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2615_update_start__ps
      -- CP-element group 134: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2615_update_start_
      -- 
    -- Element group convolve_CP_6623_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2615_update_completed__ps
      -- 
    convolve_CP_6623_elements(135) <= convolve_CP_6623_elements(136);
    -- CP-element group 136:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	135 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/type_cast_2615_update_completed_
      -- 
    -- Element group convolve_CP_6623_elements(136) is a control-delay.
    cp_element_136_delay: control_delay_element  generic map(name => " 136_delay", delay_value => 1)  port map(req => convolve_CP_6623_elements(134), ack => convolve_CP_6623_elements(136), clk => clk, reset =>reset);
    -- CP-element group 137:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (4) 
      -- CP-element group 137: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_sample_start__ps
      -- CP-element group 137: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_Sample/req
      -- 
    req_7003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(137), ack => n_chl_2951_2616_buf_req_0); -- 
    -- Element group convolve_CP_6623_elements(137) is bound as output of CP function.
    -- CP-element group 138:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_update_start__ps
      -- CP-element group 138: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_update_start_
      -- CP-element group 138: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_Update/req
      -- 
    req_7008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(138), ack => n_chl_2951_2616_buf_req_1); -- 
    -- Element group convolve_CP_6623_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (4) 
      -- CP-element group 139: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_sample_completed__ps
      -- CP-element group 139: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_Sample/ack
      -- 
    ack_7004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_2951_2616_buf_ack_0, ack => convolve_CP_6623_elements(139)); -- 
    -- CP-element group 140:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_update_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/R_n_chl_2616_Update/ack
      -- 
    ack_7009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_2951_2616_buf_ack_1, ack => convolve_CP_6623_elements(140)); -- 
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	23 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	144 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_Sample/rr
      -- 
    rr_7018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(141), ack => RPIPE_input_pipe1_2629_inst_req_0); -- 
    convolve_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(144);
      gj_convolve_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	26 
    -- CP-element group 142: 	89 
    -- CP-element group 142: 	108 
    -- CP-element group 142: 	143 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	194 
    -- CP-element group 142: 	300 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	85 
    -- CP-element group 142: 	104 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_update_start_
      -- CP-element group 142: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_Update/cr
      -- 
    cr_7023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(142), ack => RPIPE_input_pipe1_2629_inst_req_1); -- 
    convolve_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(143) & convolve_CP_6623_elements(194) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	142 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_Sample/ra
      -- 
    ra_7019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_2629_inst_ack_0, ack => convolve_CP_6623_elements(143)); -- 
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	193 
    -- CP-element group 144: 	298 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	29 
    -- CP-element group 144: 	141 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe1_2629_Update/ca
      -- 
    ca_7024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_2629_inst_ack_1, ack => convolve_CP_6623_elements(144)); -- 
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	23 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	148 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_Sample/rr
      -- 
    rr_7032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(145), ack => RPIPE_input_pipe2_2633_inst_req_0); -- 
    convolve_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(148);
      gj_convolve_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	26 
    -- CP-element group 146: 	89 
    -- CP-element group 146: 	108 
    -- CP-element group 146: 	147 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	201 
    -- CP-element group 146: 	300 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	85 
    -- CP-element group 146: 	104 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_update_start_
      -- CP-element group 146: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_Update/cr
      -- 
    cr_7037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(146), ack => RPIPE_input_pipe2_2633_inst_req_1); -- 
    convolve_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(147) & convolve_CP_6623_elements(201) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	146 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_Sample/ra
      -- 
    ra_7033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_2633_inst_ack_0, ack => convolve_CP_6623_elements(147)); -- 
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	200 
    -- CP-element group 148: 	298 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	29 
    -- CP-element group 148: 	46 
    -- CP-element group 148: 	145 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe2_2633_Update/ca
      -- 
    ca_7038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_2633_inst_ack_1, ack => convolve_CP_6623_elements(148)); -- 
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	23 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	152 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_Sample/rr
      -- 
    rr_7046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(149), ack => RPIPE_input_pipe3_2637_inst_req_0); -- 
    convolve_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(152);
      gj_convolve_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	26 
    -- CP-element group 150: 	89 
    -- CP-element group 150: 	108 
    -- CP-element group 150: 	151 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	208 
    -- CP-element group 150: 	300 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	85 
    -- CP-element group 150: 	104 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_update_start_
      -- CP-element group 150: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_Update/cr
      -- 
    cr_7051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(150), ack => RPIPE_input_pipe3_2637_inst_req_1); -- 
    convolve_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(151) & convolve_CP_6623_elements(208) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	150 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_Sample/ra
      -- 
    ra_7047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_2637_inst_ack_0, ack => convolve_CP_6623_elements(151)); -- 
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	207 
    -- CP-element group 152: 	298 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	29 
    -- CP-element group 152: 	46 
    -- CP-element group 152: 	149 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe3_2637_Update/ca
      -- 
    ca_7052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_2637_inst_ack_1, ack => convolve_CP_6623_elements(152)); -- 
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	23 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	156 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_Sample/rr
      -- 
    rr_7060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(153), ack => RPIPE_input_pipe4_2641_inst_req_0); -- 
    convolve_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(156);
      gj_convolve_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	26 
    -- CP-element group 154: 	89 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	108 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	215 
    -- CP-element group 154: 	300 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	85 
    -- CP-element group 154: 	104 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_update_start_
      -- CP-element group 154: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_Update/cr
      -- 
    cr_7065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(154), ack => RPIPE_input_pipe4_2641_inst_req_1); -- 
    convolve_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(155) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(215) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	154 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_Sample/ra
      -- 
    ra_7061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe4_2641_inst_ack_0, ack => convolve_CP_6623_elements(155)); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	214 
    -- CP-element group 156: 	298 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	46 
    -- CP-element group 156: 	153 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_input_pipe4_2641_Update/ca
      -- 
    ca_7066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe4_2641_inst_ack_1, ack => convolve_CP_6623_elements(156)); -- 
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	23 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	160 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_Sample/rr
      -- 
    rr_7074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(157), ack => RPIPE_xxconvolvexxconv_ip1_2645_inst_req_0); -- 
    convolve_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(160);
      gj_convolve_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	26 
    -- CP-element group 158: 	89 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	108 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	194 
    -- CP-element group 158: 	300 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	85 
    -- CP-element group 158: 	104 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_update_start_
      -- CP-element group 158: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_Update/cr
      -- 
    cr_7079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(158), ack => RPIPE_xxconvolvexxconv_ip1_2645_inst_req_1); -- 
    convolve_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(159) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(194) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	158 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_Sample/ra
      -- 
    ra_7075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_2645_inst_ack_0, ack => convolve_CP_6623_elements(159)); -- 
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	193 
    -- CP-element group 160: 	298 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	29 
    -- CP-element group 160: 	157 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip1_2645_Update/ca
      -- 
    ca_7080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_2645_inst_ack_1, ack => convolve_CP_6623_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	23 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	164 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_Sample/rr
      -- 
    rr_7088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(161), ack => RPIPE_xxconvolvexxconv_ip2_2649_inst_req_0); -- 
    convolve_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(164);
      gj_convolve_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	26 
    -- CP-element group 162: 	89 
    -- CP-element group 162: 	108 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	201 
    -- CP-element group 162: 	300 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	85 
    -- CP-element group 162: 	104 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_update_start_
      -- CP-element group 162: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_Update/cr
      -- 
    cr_7093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(162), ack => RPIPE_xxconvolvexxconv_ip2_2649_inst_req_1); -- 
    convolve_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(163) & convolve_CP_6623_elements(26) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(201) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	162 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_Sample/ra
      -- 
    ra_7089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_2649_inst_ack_0, ack => convolve_CP_6623_elements(163)); -- 
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	200 
    -- CP-element group 164: 	298 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	161 
    -- CP-element group 164: 	29 
    -- CP-element group 164: 	46 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip2_2649_Update/ca
      -- 
    ca_7094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_2649_inst_ack_1, ack => convolve_CP_6623_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	23 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	168 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_Sample/rr
      -- 
    rr_7102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(165), ack => RPIPE_xxconvolvexxconv_ip3_2653_inst_req_0); -- 
    convolve_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(168);
      gj_convolve_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	26 
    -- CP-element group 166: 	89 
    -- CP-element group 166: 	167 
    -- CP-element group 166: 	108 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	208 
    -- CP-element group 166: 	300 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	85 
    -- CP-element group 166: 	104 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_update_start_
      -- CP-element group 166: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_Update/cr
      -- 
    cr_7107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(166), ack => RPIPE_xxconvolvexxconv_ip3_2653_inst_req_1); -- 
    convolve_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(167) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(208) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	166 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_Sample/ra
      -- 
    ra_7103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_2653_inst_ack_0, ack => convolve_CP_6623_elements(167)); -- 
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	207 
    -- CP-element group 168: 	298 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	165 
    -- CP-element group 168: 	29 
    -- CP-element group 168: 	46 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip3_2653_Update/ca
      -- 
    ca_7108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_2653_inst_ack_1, ack => convolve_CP_6623_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	23 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	172 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_Sample/rr
      -- 
    rr_7116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(169), ack => RPIPE_xxconvolvexxconv_ip4_2657_inst_req_0); -- 
    convolve_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(172);
      gj_convolve_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	26 
    -- CP-element group 170: 	89 
    -- CP-element group 170: 	171 
    -- CP-element group 170: 	108 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	215 
    -- CP-element group 170: 	300 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	85 
    -- CP-element group 170: 	104 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_update_start_
      -- CP-element group 170: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_Update/cr
      -- 
    cr_7121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(170), ack => RPIPE_xxconvolvexxconv_ip4_2657_inst_req_1); -- 
    convolve_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(171) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(215) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	170 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_Sample/ra
      -- 
    ra_7117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip4_2657_inst_ack_0, ack => convolve_CP_6623_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	214 
    -- CP-element group 172: 	298 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	46 
    -- CP-element group 172: 	169 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_ip4_2657_Update/ca
      -- 
    ca_7122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip4_2657_inst_ack_1, ack => convolve_CP_6623_elements(172)); -- 
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	89 
    -- CP-element group 173: 	108 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_Sample/req
      -- 
    req_7130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(173), ack => W_read_ip_2603_delayed_1_0_2659_inst_req_0); -- 
    convolve_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(175);
      gj_convolve_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	26 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	194 
    -- CP-element group 174: 	176 
    -- CP-element group 174: 	300 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_update_start_
      -- CP-element group 174: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_Update/req
      -- 
    req_7135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(174), ack => W_read_ip_2603_delayed_1_0_2659_inst_req_1); -- 
    convolve_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(194) & convolve_CP_6623_elements(176) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	85 
    -- CP-element group 175: 	173 
    -- CP-element group 175: 	104 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_Sample/ack
      -- 
    ack_7131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2603_delayed_1_0_2659_inst_ack_0, ack => convolve_CP_6623_elements(175)); -- 
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	193 
    -- CP-element group 176: 	298 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	29 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2661_Update/ack
      -- 
    ack_7136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2603_delayed_1_0_2659_inst_ack_1, ack => convolve_CP_6623_elements(176)); -- 
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	89 
    -- CP-element group 177: 	108 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_Sample/req
      -- 
    req_7144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(177), ack => W_read_ip_2609_delayed_1_0_2668_inst_req_0); -- 
    convolve_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(179);
      gj_convolve_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	26 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	201 
    -- CP-element group 178: 	180 
    -- CP-element group 178: 	300 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_update_start_
      -- CP-element group 178: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_Update/req
      -- 
    req_7149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(178), ack => W_read_ip_2609_delayed_1_0_2668_inst_req_1); -- 
    convolve_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(201) & convolve_CP_6623_elements(180) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	85 
    -- CP-element group 179: 	104 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_Sample/ack
      -- 
    ack_7145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2609_delayed_1_0_2668_inst_ack_0, ack => convolve_CP_6623_elements(179)); -- 
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	200 
    -- CP-element group 180: 	298 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	29 
    -- CP-element group 180: 	46 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2670_Update/ack
      -- 
    ack_7150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2609_delayed_1_0_2668_inst_ack_1, ack => convolve_CP_6623_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	89 
    -- CP-element group 181: 	108 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_Sample/req
      -- 
    req_7158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(181), ack => W_read_ip_2615_delayed_1_0_2677_inst_req_0); -- 
    convolve_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(183);
      gj_convolve_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	26 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: 	208 
    -- CP-element group 182: 	300 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_update_start_
      -- CP-element group 182: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_Update/req
      -- 
    req_7163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(182), ack => W_read_ip_2615_delayed_1_0_2677_inst_req_1); -- 
    convolve_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(184) & convolve_CP_6623_elements(208) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	85 
    -- CP-element group 183: 	181 
    -- CP-element group 183: 	104 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_Sample/ack
      -- 
    ack_7159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2615_delayed_1_0_2677_inst_ack_0, ack => convolve_CP_6623_elements(183)); -- 
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	207 
    -- CP-element group 184: 	298 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	29 
    -- CP-element group 184: 	46 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2679_Update/ack
      -- 
    ack_7164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2615_delayed_1_0_2677_inst_ack_1, ack => convolve_CP_6623_elements(184)); -- 
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	89 
    -- CP-element group 185: 	108 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_Sample/req
      -- 
    req_7172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(185), ack => W_read_ip_2621_delayed_1_0_2686_inst_req_0); -- 
    convolve_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(187);
      gj_convolve_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	26 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	215 
    -- CP-element group 186: 	188 
    -- CP-element group 186: 	300 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_update_start_
      -- CP-element group 186: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_Update/req
      -- 
    req_7177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(186), ack => W_read_ip_2621_delayed_1_0_2686_inst_req_1); -- 
    convolve_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(215) & convolve_CP_6623_elements(188) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	85 
    -- CP-element group 187: 	185 
    -- CP-element group 187: 	104 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_Sample/ack
      -- 
    ack_7173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2621_delayed_1_0_2686_inst_ack_0, ack => convolve_CP_6623_elements(187)); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	214 
    -- CP-element group 188: 	298 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	46 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2688_Update/ack
      -- 
    ack_7178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2621_delayed_1_0_2686_inst_ack_1, ack => convolve_CP_6623_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	89 
    -- CP-element group 189: 	108 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_Sample/req
      -- 
    req_7186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(189), ack => W_write_input_2635_delayed_1_0_2704_inst_req_0); -- 
    convolve_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(191);
      gj_convolve_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_update_start_
      -- CP-element group 190: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_Update/req
      -- 
    req_7191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(190), ack => W_write_input_2635_delayed_1_0_2704_inst_req_1); -- 
    convolve_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(194) & convolve_CP_6623_elements(192);
      gj_convolve_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	85 
    -- CP-element group 191: 	189 
    -- CP-element group 191: 	104 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_Sample/ack
      -- 
    ack_7187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2635_delayed_1_0_2704_inst_ack_0, ack => convolve_CP_6623_elements(191)); -- 
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2706_Update/ack
      -- 
    ack_7192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2635_delayed_1_0_2704_inst_ack_1, ack => convolve_CP_6623_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	160 
    -- CP-element group 193: 	192 
    -- CP-element group 193: 	144 
    -- CP-element group 193: 	176 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_Sample/req
      -- 
    req_7200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(193), ack => WPIPE_xxconvolvexxconv_ip1_2708_inst_req_0); -- 
    convolve_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(160) & convolve_CP_6623_elements(192) & convolve_CP_6623_elements(144) & convolve_CP_6623_elements(176) & convolve_CP_6623_elements(195);
      gj_convolve_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	158 
    -- CP-element group 194: 	190 
    -- CP-element group 194: 	142 
    -- CP-element group 194: 	174 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_update_start_
      -- CP-element group 194: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_Update/req
      -- 
    ack_7201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_2708_inst_ack_0, ack => convolve_CP_6623_elements(194)); -- 
    req_7205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(194), ack => WPIPE_xxconvolvexxconv_ip1_2708_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	306 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip1_2708_Update/ack
      -- 
    ack_7206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_2708_inst_ack_1, ack => convolve_CP_6623_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	89 
    -- CP-element group 196: 	108 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_Sample/req
      -- 
    req_7214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(196), ack => W_write_input_2639_delayed_1_0_2711_inst_req_0); -- 
    convolve_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(198);
      gj_convolve_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	199 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_update_start_
      -- CP-element group 197: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_Update/req
      -- 
    req_7219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(197), ack => W_write_input_2639_delayed_1_0_2711_inst_req_1); -- 
    convolve_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(199) & convolve_CP_6623_elements(201);
      gj_convolve_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: 	85 
    -- CP-element group 198: 	104 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_Sample/ack
      -- 
    ack_7215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2639_delayed_1_0_2711_inst_ack_0, ack => convolve_CP_6623_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	197 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2713_Update/ack
      -- 
    ack_7220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2639_delayed_1_0_2711_inst_ack_1, ack => convolve_CP_6623_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	164 
    -- CP-element group 200: 	199 
    -- CP-element group 200: 	180 
    -- CP-element group 200: 	148 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_Sample/req
      -- 
    req_7228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(200), ack => WPIPE_xxconvolvexxconv_ip2_2715_inst_req_0); -- 
    convolve_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(164) & convolve_CP_6623_elements(199) & convolve_CP_6623_elements(180) & convolve_CP_6623_elements(148) & convolve_CP_6623_elements(202);
      gj_convolve_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	197 
    -- CP-element group 201: 	162 
    -- CP-element group 201: 	146 
    -- CP-element group 201: 	178 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_update_start_
      -- CP-element group 201: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_Update/req
      -- 
    ack_7229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_2715_inst_ack_0, ack => convolve_CP_6623_elements(201)); -- 
    req_7233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(201), ack => WPIPE_xxconvolvexxconv_ip2_2715_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	306 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip2_2715_Update/ack
      -- 
    ack_7234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_2715_inst_ack_1, ack => convolve_CP_6623_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	89 
    -- CP-element group 203: 	108 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	205 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_Sample/req
      -- 
    req_7242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(203), ack => W_write_input_2643_delayed_1_0_2718_inst_req_0); -- 
    convolve_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(205);
      gj_convolve_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	206 
    -- CP-element group 204: 	208 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_update_start_
      -- CP-element group 204: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_Update/req
      -- 
    req_7247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(204), ack => W_write_input_2643_delayed_1_0_2718_inst_req_1); -- 
    convolve_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(206) & convolve_CP_6623_elements(208);
      gj_convolve_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	85 
    -- CP-element group 205: 	203 
    -- CP-element group 205: 	104 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_Sample/ack
      -- 
    ack_7243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2643_delayed_1_0_2718_inst_ack_0, ack => convolve_CP_6623_elements(205)); -- 
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2720_Update/ack
      -- 
    ack_7248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2643_delayed_1_0_2718_inst_ack_1, ack => convolve_CP_6623_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	168 
    -- CP-element group 207: 	184 
    -- CP-element group 207: 	152 
    -- CP-element group 207: 	206 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_Sample/req
      -- 
    req_7256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(207), ack => WPIPE_xxconvolvexxconv_ip3_2722_inst_req_0); -- 
    convolve_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(168) & convolve_CP_6623_elements(184) & convolve_CP_6623_elements(152) & convolve_CP_6623_elements(206) & convolve_CP_6623_elements(209);
      gj_convolve_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	166 
    -- CP-element group 208: 	204 
    -- CP-element group 208: 	182 
    -- CP-element group 208: 	150 
    -- CP-element group 208:  members (6) 
      -- CP-element group 208: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_update_start_
      -- CP-element group 208: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_Sample/ack
      -- CP-element group 208: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_Update/req
      -- 
    ack_7257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_2722_inst_ack_0, ack => convolve_CP_6623_elements(208)); -- 
    req_7261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(208), ack => WPIPE_xxconvolvexxconv_ip3_2722_inst_req_1); -- 
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	306 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	207 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip3_2722_Update/ack
      -- 
    ack_7262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_2722_inst_ack_1, ack => convolve_CP_6623_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	89 
    -- CP-element group 210: 	108 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_Sample/req
      -- 
    req_7270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(210), ack => W_write_input_2647_delayed_1_0_2725_inst_req_0); -- 
    convolve_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(89) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(212);
      gj_convolve_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: 	215 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_update_start_
      -- CP-element group 211: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_Update/req
      -- 
    req_7275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(211), ack => W_write_input_2647_delayed_1_0_2725_inst_req_1); -- 
    convolve_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(213) & convolve_CP_6623_elements(215);
      gj_convolve_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: 	85 
    -- CP-element group 212: 	104 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_Sample/ack
      -- 
    ack_7271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2647_delayed_1_0_2725_inst_ack_0, ack => convolve_CP_6623_elements(212)); -- 
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2727_Update/ack
      -- 
    ack_7276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2647_delayed_1_0_2725_inst_ack_1, ack => convolve_CP_6623_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: 	172 
    -- CP-element group 214: 	156 
    -- CP-element group 214: 	188 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_Sample/req
      -- 
    req_7284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(214), ack => WPIPE_xxconvolvexxconv_ip4_2729_inst_req_0); -- 
    convolve_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(213) & convolve_CP_6623_elements(172) & convolve_CP_6623_elements(156) & convolve_CP_6623_elements(188) & convolve_CP_6623_elements(216);
      gj_convolve_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	211 
    -- CP-element group 215: 	170 
    -- CP-element group 215: 	154 
    -- CP-element group 215: 	186 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_update_start_
      -- CP-element group 215: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_Sample/ack
      -- CP-element group 215: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_Update/req
      -- 
    ack_7285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip4_2729_inst_ack_0, ack => convolve_CP_6623_elements(215)); -- 
    req_7289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(215), ack => WPIPE_xxconvolvexxconv_ip4_2729_inst_req_1); -- 
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	306 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_ip4_2729_Update/ack
      -- 
    ack_7290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip4_2729_inst_ack_1, ack => convolve_CP_6623_elements(216)); -- 
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	23 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	220 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_sample_start_
      -- CP-element group 217: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_Sample/$entry
      -- CP-element group 217: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_Sample/rr
      -- 
    rr_7298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(217), ack => RPIPE_kernel_pipe1_2759_inst_req_0); -- 
    convolve_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(220);
      gj_convolve_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	219 
    -- CP-element group 218: 	26 
    -- CP-element group 218: 	70 
    -- CP-element group 218: 	89 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	270 
    -- CP-element group 218: 	300 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	66 
    -- CP-element group 218: 	85 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_update_start_
      -- CP-element group 218: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_Update/cr
      -- 
    cr_7303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(218), ack => RPIPE_kernel_pipe1_2759_inst_req_1); -- 
    convolve_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(219) & convolve_CP_6623_elements(26) & convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(270) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	218 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_Sample/ra
      -- 
    ra_7299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_2759_inst_ack_0, ack => convolve_CP_6623_elements(219)); -- 
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	269 
    -- CP-element group 220: 	298 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	217 
    -- CP-element group 220: 	29 
    -- CP-element group 220: 	46 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe1_2759_Update/ca
      -- 
    ca_7304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_2759_inst_ack_1, ack => convolve_CP_6623_elements(220)); -- 
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	23 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	224 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_sample_start_
      -- CP-element group 221: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_Sample/rr
      -- 
    rr_7312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(221), ack => RPIPE_kernel_pipe2_2763_inst_req_0); -- 
    convolve_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(224);
      gj_convolve_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	223 
    -- CP-element group 222: 	26 
    -- CP-element group 222: 	70 
    -- CP-element group 222: 	89 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	277 
    -- CP-element group 222: 	300 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	66 
    -- CP-element group 222: 	85 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_update_start_
      -- CP-element group 222: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_Update/$entry
      -- CP-element group 222: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_Update/cr
      -- 
    cr_7317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(222), ack => RPIPE_kernel_pipe2_2763_inst_req_1); -- 
    convolve_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(223) & convolve_CP_6623_elements(26) & convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(277) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	222 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_Sample/ra
      -- 
    ra_7313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_2763_inst_ack_0, ack => convolve_CP_6623_elements(223)); -- 
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	276 
    -- CP-element group 224: 	298 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	221 
    -- CP-element group 224: 	29 
    -- CP-element group 224: 	46 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe2_2763_Update/ca
      -- 
    ca_7318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_2763_inst_ack_1, ack => convolve_CP_6623_elements(224)); -- 
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	23 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	228 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_Sample/rr
      -- 
    rr_7326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(225), ack => RPIPE_kernel_pipe3_2767_inst_req_0); -- 
    convolve_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(228);
      gj_convolve_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	227 
    -- CP-element group 226: 	26 
    -- CP-element group 226: 	70 
    -- CP-element group 226: 	89 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	284 
    -- CP-element group 226: 	300 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: marked-successors 
    -- CP-element group 226: 	66 
    -- CP-element group 226: 	85 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_update_start_
      -- CP-element group 226: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_Update/cr
      -- 
    cr_7331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(226), ack => RPIPE_kernel_pipe3_2767_inst_req_1); -- 
    convolve_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(227) & convolve_CP_6623_elements(26) & convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(284) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	226 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_Sample/ra
      -- 
    ra_7327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_2767_inst_ack_0, ack => convolve_CP_6623_elements(227)); -- 
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	283 
    -- CP-element group 228: 	298 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	225 
    -- CP-element group 228: 	29 
    -- CP-element group 228: 	46 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_kernel_pipe3_2767_Update/ca
      -- 
    ca_7332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_2767_inst_ack_1, ack => convolve_CP_6623_elements(228)); -- 
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	23 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	232 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_Sample/rr
      -- 
    rr_7340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(229), ack => RPIPE_xxconvolvexxconv_k1_2771_inst_req_0); -- 
    convolve_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(232);
      gj_convolve_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	231 
    -- CP-element group 230: 	26 
    -- CP-element group 230: 	70 
    -- CP-element group 230: 	89 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	270 
    -- CP-element group 230: 	300 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	66 
    -- CP-element group 230: 	85 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_update_start_
      -- CP-element group 230: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_Update/cr
      -- 
    cr_7345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(230), ack => RPIPE_xxconvolvexxconv_k1_2771_inst_req_1); -- 
    convolve_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(231) & convolve_CP_6623_elements(26) & convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(270) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	230 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_Sample/ra
      -- 
    ra_7341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_2771_inst_ack_0, ack => convolve_CP_6623_elements(231)); -- 
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	269 
    -- CP-element group 232: 	298 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	229 
    -- CP-element group 232: 	29 
    -- CP-element group 232: 	46 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k1_2771_Update/ca
      -- 
    ca_7346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_2771_inst_ack_1, ack => convolve_CP_6623_elements(232)); -- 
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	23 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	236 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_Sample/rr
      -- 
    rr_7354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(233), ack => RPIPE_xxconvolvexxconv_k2_2775_inst_req_0); -- 
    convolve_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(236);
      gj_convolve_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	26 
    -- CP-element group 234: 	70 
    -- CP-element group 234: 	89 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	277 
    -- CP-element group 234: 	300 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: marked-successors 
    -- CP-element group 234: 	66 
    -- CP-element group 234: 	85 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_update_start_
      -- CP-element group 234: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_Update/cr
      -- 
    cr_7359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(234), ack => RPIPE_xxconvolvexxconv_k2_2775_inst_req_1); -- 
    convolve_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(235) & convolve_CP_6623_elements(26) & convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(277) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	234 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_Sample/ra
      -- 
    ra_7355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_2775_inst_ack_0, ack => convolve_CP_6623_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	276 
    -- CP-element group 236: 	298 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	233 
    -- CP-element group 236: 	29 
    -- CP-element group 236: 	46 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k2_2775_Update/ca
      -- 
    ca_7360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_2775_inst_ack_1, ack => convolve_CP_6623_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	23 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	240 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_Sample/rr
      -- 
    rr_7368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(237), ack => RPIPE_xxconvolvexxconv_k3_2779_inst_req_0); -- 
    convolve_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(240);
      gj_convolve_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	239 
    -- CP-element group 238: 	26 
    -- CP-element group 238: 	70 
    -- CP-element group 238: 	89 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	284 
    -- CP-element group 238: 	300 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	66 
    -- CP-element group 238: 	85 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_update_start_
      -- CP-element group 238: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_Update/cr
      -- 
    cr_7373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(238), ack => RPIPE_xxconvolvexxconv_k3_2779_inst_req_1); -- 
    convolve_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(239) & convolve_CP_6623_elements(26) & convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(284) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	238 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_Sample/ra
      -- 
    ra_7369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_2779_inst_ack_0, ack => convolve_CP_6623_elements(239)); -- 
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	283 
    -- CP-element group 240: 	298 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	237 
    -- CP-element group 240: 	29 
    -- CP-element group 240: 	46 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/RPIPE_xxconvolvexxconv_k3_2779_Update/ca
      -- 
    ca_7374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_2779_inst_ack_1, ack => convolve_CP_6623_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	70 
    -- CP-element group 241: 	89 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_Sample/req
      -- 
    req_7382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(241), ack => W_read_k_2701_delayed_1_0_2781_inst_req_0); -- 
    convolve_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(243);
      gj_convolve_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	26 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	244 
    -- CP-element group 242: 	270 
    -- CP-element group 242: 	300 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_update_start_
      -- CP-element group 242: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_Update/req
      -- 
    req_7387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(242), ack => W_read_k_2701_delayed_1_0_2781_inst_req_1); -- 
    convolve_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(244) & convolve_CP_6623_elements(270) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	66 
    -- CP-element group 243: 	85 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_Sample/ack
      -- 
    ack_7383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2701_delayed_1_0_2781_inst_ack_0, ack => convolve_CP_6623_elements(243)); -- 
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	269 
    -- CP-element group 244: 	298 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	29 
    -- CP-element group 244: 	46 
    -- CP-element group 244: 	242 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2783_Update/ack
      -- 
    ack_7388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2701_delayed_1_0_2781_inst_ack_1, ack => convolve_CP_6623_elements(244)); -- 
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	70 
    -- CP-element group 245: 	89 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_Sample/req
      -- 
    req_7396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(245), ack => W_read_k_2707_delayed_1_0_2790_inst_req_0); -- 
    convolve_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(247);
      gj_convolve_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	26 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	248 
    -- CP-element group 246: 	277 
    -- CP-element group 246: 	300 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_update_start_
      -- CP-element group 246: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_Update/req
      -- 
    req_7401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(246), ack => W_read_k_2707_delayed_1_0_2790_inst_req_1); -- 
    convolve_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(248) & convolve_CP_6623_elements(277) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	66 
    -- CP-element group 247: 	85 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_Sample/ack
      -- 
    ack_7397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2707_delayed_1_0_2790_inst_ack_0, ack => convolve_CP_6623_elements(247)); -- 
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	276 
    -- CP-element group 248: 	298 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	29 
    -- CP-element group 248: 	46 
    -- CP-element group 248: 	246 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2792_Update/ack
      -- 
    ack_7402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2707_delayed_1_0_2790_inst_ack_1, ack => convolve_CP_6623_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	70 
    -- CP-element group 249: 	89 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_Sample/req
      -- 
    req_7410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(249), ack => W_read_k_2713_delayed_1_0_2799_inst_req_0); -- 
    convolve_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(251);
      gj_convolve_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	26 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	252 
    -- CP-element group 250: 	284 
    -- CP-element group 250: 	300 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_update_start_
      -- CP-element group 250: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_Update/req
      -- 
    req_7415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(250), ack => W_read_k_2713_delayed_1_0_2799_inst_req_1); -- 
    convolve_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(252) & convolve_CP_6623_elements(284) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	66 
    -- CP-element group 251: 	85 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_Sample/ack
      -- 
    ack_7411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2713_delayed_1_0_2799_inst_ack_0, ack => convolve_CP_6623_elements(251)); -- 
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	283 
    -- CP-element group 252: 	298 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	29 
    -- CP-element group 252: 	46 
    -- CP-element group 252: 	250 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2801_Update/ack
      -- 
    ack_7416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2713_delayed_1_0_2799_inst_ack_1, ack => convolve_CP_6623_elements(252)); -- 
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	32 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_Sample/req
      -- 
    req_7424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(253), ack => W_acc1_2767_delayed_1_0_2856_inst_req_0); -- 
    convolve_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(32) & convolve_CP_6623_elements(255);
      gj_convolve_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	26 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: 	300 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_update_start_
      -- CP-element group 254: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_Update/req
      -- 
    req_7429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(254), ack => W_acc1_2767_delayed_1_0_2856_inst_req_1); -- 
    convolve_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(256) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	30 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_Sample/ack
      -- 
    ack_7425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc1_2767_delayed_1_0_2856_inst_ack_0, ack => convolve_CP_6623_elements(255)); -- 
    -- CP-element group 256:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	298 
    -- CP-element group 256: marked-successors 
    -- CP-element group 256: 	29 
    -- CP-element group 256: 	254 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2858_Update/ack
      -- 
    ack_7430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc1_2767_delayed_1_0_2856_inst_ack_1, ack => convolve_CP_6623_elements(256)); -- 
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	51 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_sample_start_
      -- CP-element group 257: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_Sample/$entry
      -- CP-element group 257: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_Sample/req
      -- 
    req_7438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(257), ack => W_acc2_2776_delayed_1_0_2868_inst_req_0); -- 
    convolve_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(51) & convolve_CP_6623_elements(259);
      gj_convolve_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	26 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: 	300 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_update_start_
      -- CP-element group 258: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_Update/req
      -- 
    req_7443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(258), ack => W_acc2_2776_delayed_1_0_2868_inst_req_1); -- 
    convolve_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(260) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	47 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_sample_completed_
      -- CP-element group 259: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_Sample/ack
      -- 
    ack_7439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc2_2776_delayed_1_0_2868_inst_ack_0, ack => convolve_CP_6623_elements(259)); -- 
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	298 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	46 
    -- CP-element group 260: 	258 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2870_Update/ack
      -- 
    ack_7444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc2_2776_delayed_1_0_2868_inst_ack_1, ack => convolve_CP_6623_elements(260)); -- 
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	23 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_Sample/rr
      -- 
    rr_7452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(261), ack => SUB_u16_u16_2905_inst_req_0); -- 
    convolve_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(23) & convolve_CP_6623_elements(263);
      gj_convolve_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	264 
    -- CP-element group 262: 	267 
    -- CP-element group 262: 	274 
    -- CP-element group 262: 	281 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_update_start_
      -- CP-element group 262: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_Update/$entry
      -- 
    cr_7457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(262), ack => SUB_u16_u16_2905_inst_req_1); -- 
    convolve_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(264) & convolve_CP_6623_elements(267) & convolve_CP_6623_elements(274) & convolve_CP_6623_elements(281);
      gj_convolve_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_Sample/ra
      -- 
    ra_7453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2905_inst_ack_0, ack => convolve_CP_6623_elements(263)); -- 
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	24 
    -- CP-element group 264: 	265 
    -- CP-element group 264: 	272 
    -- CP-element group 264: 	279 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/SUB_u16_u16_2905_Update/ca
      -- 
    ca_7458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2905_inst_ack_1, ack => convolve_CP_6623_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	70 
    -- CP-element group 265: 	89 
    -- CP-element group 265: 	264 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_Sample/req
      -- CP-element group 265: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_Sample/$entry
      -- 
    req_7466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(265), ack => W_store_kernel_2824_delayed_1_0_2923_inst_req_0); -- 
    convolve_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(264) & convolve_CP_6623_elements(267);
      gj_convolve_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: 	270 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_Update/req
      -- CP-element group 266: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_update_start_
      -- 
    req_7471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(266), ack => W_store_kernel_2824_delayed_1_0_2923_inst_req_1); -- 
    convolve_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(268) & convolve_CP_6623_elements(270);
      gj_convolve_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	66 
    -- CP-element group 267: 	85 
    -- CP-element group 267: 	262 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_Sample/ack
      -- 
    ack_7467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2824_delayed_1_0_2923_inst_ack_0, ack => convolve_CP_6623_elements(267)); -- 
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2925_update_completed_
      -- 
    ack_7472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2824_delayed_1_0_2923_inst_ack_1, ack => convolve_CP_6623_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	232 
    -- CP-element group 269: 	220 
    -- CP-element group 269: 	244 
    -- CP-element group 269: 	268 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_Sample/req
      -- CP-element group 269: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_sample_start_
      -- 
    req_7480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(269), ack => WPIPE_xxconvolvexxconv_k1_2927_inst_req_0); -- 
    convolve_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(232) & convolve_CP_6623_elements(220) & convolve_CP_6623_elements(244) & convolve_CP_6623_elements(268) & convolve_CP_6623_elements(271);
      gj_convolve_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	230 
    -- CP-element group 270: 	218 
    -- CP-element group 270: 	242 
    -- CP-element group 270: 	266 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_update_start_
      -- CP-element group 270: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_Sample/ack
      -- CP-element group 270: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_Update/req
      -- 
    ack_7481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_2927_inst_ack_0, ack => convolve_CP_6623_elements(270)); -- 
    req_7485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(270), ack => WPIPE_xxconvolvexxconv_k1_2927_inst_req_1); -- 
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	306 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k1_2927_Update/ack
      -- 
    ack_7486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_2927_inst_ack_1, ack => convolve_CP_6623_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	70 
    -- CP-element group 272: 	89 
    -- CP-element group 272: 	264 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_Sample/req
      -- 
    req_7494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(272), ack => W_store_kernel_2828_delayed_1_0_2930_inst_req_0); -- 
    convolve_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(264) & convolve_CP_6623_elements(274);
      gj_convolve_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: 	277 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_update_start_
      -- CP-element group 273: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_Update/req
      -- 
    req_7499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(273), ack => W_store_kernel_2828_delayed_1_0_2930_inst_req_1); -- 
    convolve_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(275) & convolve_CP_6623_elements(277);
      gj_convolve_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	66 
    -- CP-element group 274: 	85 
    -- CP-element group 274: 	262 
    -- CP-element group 274: 	272 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_Sample/ack
      -- CP-element group 274: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_sample_completed_
      -- 
    ack_7495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2828_delayed_1_0_2930_inst_ack_0, ack => convolve_CP_6623_elements(274)); -- 
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_update_completed_
      -- CP-element group 275: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2932_Update/ack
      -- 
    ack_7500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2828_delayed_1_0_2930_inst_ack_1, ack => convolve_CP_6623_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	224 
    -- CP-element group 276: 	236 
    -- CP-element group 276: 	248 
    -- CP-element group 276: 	275 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_sample_start_
      -- 
    req_7508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(276), ack => WPIPE_xxconvolvexxconv_k2_2934_inst_req_0); -- 
    convolve_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(224) & convolve_CP_6623_elements(236) & convolve_CP_6623_elements(248) & convolve_CP_6623_elements(275) & convolve_CP_6623_elements(278);
      gj_convolve_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277: marked-successors 
    -- CP-element group 277: 	234 
    -- CP-element group 277: 	222 
    -- CP-element group 277: 	246 
    -- CP-element group 277: 	273 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_update_start_
      -- CP-element group 277: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_Update/req
      -- CP-element group 277: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_sample_completed_
      -- 
    ack_7509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_2934_inst_ack_0, ack => convolve_CP_6623_elements(277)); -- 
    req_7513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(277), ack => WPIPE_xxconvolvexxconv_k2_2934_inst_req_1); -- 
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	306 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k2_2934_Update/$exit
      -- 
    ack_7514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_2934_inst_ack_1, ack => convolve_CP_6623_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	70 
    -- CP-element group 279: 	89 
    -- CP-element group 279: 	264 
    -- CP-element group 279: marked-predecessors 
    -- CP-element group 279: 	281 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_Sample/req
      -- CP-element group 279: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_sample_start_
      -- 
    req_7522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(279), ack => W_store_kernel_2832_delayed_1_0_2937_inst_req_0); -- 
    convolve_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(70) & convolve_CP_6623_elements(89) & convolve_CP_6623_elements(264) & convolve_CP_6623_elements(281);
      gj_convolve_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: marked-predecessors 
    -- CP-element group 280: 	282 
    -- CP-element group 280: 	284 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_update_start_
      -- CP-element group 280: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_Update/req
      -- CP-element group 280: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_Update/$entry
      -- 
    req_7527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(280), ack => W_store_kernel_2832_delayed_1_0_2937_inst_req_1); -- 
    convolve_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(282) & convolve_CP_6623_elements(284);
      gj_convolve_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: successors 
    -- CP-element group 281: marked-successors 
    -- CP-element group 281: 	66 
    -- CP-element group 281: 	85 
    -- CP-element group 281: 	262 
    -- CP-element group 281: 	279 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_Sample/ack
      -- 
    ack_7523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2832_delayed_1_0_2937_inst_ack_0, ack => convolve_CP_6623_elements(281)); -- 
    -- CP-element group 282:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282: marked-successors 
    -- CP-element group 282: 	280 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_Update/ack
      -- CP-element group 282: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2939_Update/$exit
      -- 
    ack_7528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2832_delayed_1_0_2937_inst_ack_1, ack => convolve_CP_6623_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	228 
    -- CP-element group 283: 	240 
    -- CP-element group 283: 	252 
    -- CP-element group 283: 	282 
    -- CP-element group 283: marked-predecessors 
    -- CP-element group 283: 	285 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_Sample/$entry
      -- 
    req_7536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(283), ack => WPIPE_xxconvolvexxconv_k3_2941_inst_req_0); -- 
    convolve_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(228) & convolve_CP_6623_elements(240) & convolve_CP_6623_elements(252) & convolve_CP_6623_elements(282) & convolve_CP_6623_elements(285);
      gj_convolve_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284: marked-successors 
    -- CP-element group 284: 	226 
    -- CP-element group 284: 	238 
    -- CP-element group 284: 	250 
    -- CP-element group 284: 	280 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_Update/req
      -- CP-element group 284: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_update_start_
      -- CP-element group 284: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_Sample/$exit
      -- 
    ack_7537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_2941_inst_ack_0, ack => convolve_CP_6623_elements(284)); -- 
    req_7541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(284), ack => WPIPE_xxconvolvexxconv_k3_2941_inst_req_1); -- 
    -- CP-element group 285:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	306 
    -- CP-element group 285: marked-successors 
    -- CP-element group 285: 	283 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_Update/ack
      -- CP-element group 285: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_xxconvolvexxconv_k3_2941_update_completed_
      -- 
    ack_7542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_2941_inst_ack_1, ack => convolve_CP_6623_elements(285)); -- 
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	127 
    -- CP-element group 286: 	108 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	288 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_sample_start_
      -- CP-element group 286: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_Sample/req
      -- 
    req_7550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(286), ack => W_num_done_2875_delayed_1_0_2982_inst_req_0); -- 
    convolve_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(127) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(288);
      gj_convolve_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	26 
    -- CP-element group 287: marked-predecessors 
    -- CP-element group 287: 	289 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	289 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_Update/req
      -- CP-element group 287: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_update_start_
      -- 
    req_7555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(287), ack => W_num_done_2875_delayed_1_0_2982_inst_req_1); -- 
    convolve_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(289);
      gj_convolve_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	123 
    -- CP-element group 288: 	104 
    -- CP-element group 288: 	286 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_Sample/ack
      -- 
    ack_7551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2875_delayed_1_0_2982_inst_ack_0, ack => convolve_CP_6623_elements(288)); -- 
    -- CP-element group 289:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	287 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	306 
    -- CP-element group 289: marked-successors 
    -- CP-element group 289: 	29 
    -- CP-element group 289: 	287 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_Update/ack
      -- CP-element group 289: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2984_update_completed_
      -- 
    ack_7556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2875_delayed_1_0_2982_inst_ack_1, ack => convolve_CP_6623_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	127 
    -- CP-element group 290: 	108 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_sample_start_
      -- 
    req_7564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(290), ack => W_num_done_2881_delayed_1_0_2991_inst_req_0); -- 
    convolve_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(127) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(292);
      gj_convolve_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	26 
    -- CP-element group 291: marked-predecessors 
    -- CP-element group 291: 	293 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_update_start_
      -- CP-element group 291: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_Update/req
      -- 
    req_7569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(291), ack => W_num_done_2881_delayed_1_0_2991_inst_req_1); -- 
    convolve_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(26) & convolve_CP_6623_elements(293);
      gj_convolve_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	123 
    -- CP-element group 292: 	104 
    -- CP-element group 292: 	290 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_Sample/ack
      -- CP-element group 292: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_sample_completed_
      -- 
    ack_7565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2881_delayed_1_0_2991_inst_ack_0, ack => convolve_CP_6623_elements(292)); -- 
    -- CP-element group 293:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	306 
    -- CP-element group 293: marked-successors 
    -- CP-element group 293: 	46 
    -- CP-element group 293: 	291 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_2993_Update/ack
      -- 
    ack_7570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2881_delayed_1_0_2991_inst_ack_1, ack => convolve_CP_6623_elements(293)); -- 
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	127 
    -- CP-element group 294: 	108 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_Sample/req
      -- 
    req_7578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(294), ack => W_num_done_2886_delayed_1_0_3000_inst_req_0); -- 
    convolve_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(127) & convolve_CP_6623_elements(108) & convolve_CP_6623_elements(296);
      gj_convolve_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: marked-predecessors 
    -- CP-element group 295: 	297 
    -- CP-element group 295: 	300 
    -- CP-element group 295: 	303 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	297 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_update_start_
      -- CP-element group 295: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_Update/req
      -- 
    req_7583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(295), ack => W_num_done_2886_delayed_1_0_3000_inst_req_1); -- 
    convolve_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(297) & convolve_CP_6623_elements(300) & convolve_CP_6623_elements(303);
      gj_convolve_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	123 
    -- CP-element group 296: 	104 
    -- CP-element group 296: 	294 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_sample_completed_
      -- CP-element group 296: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_Sample/ack
      -- 
    ack_7579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2886_delayed_1_0_3000_inst_ack_0, ack => convolve_CP_6623_elements(296)); -- 
    -- CP-element group 297:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	295 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297: 	302 
    -- CP-element group 297: marked-successors 
    -- CP-element group 297: 	295 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_update_completed_
      -- CP-element group 297: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/assign_stmt_3002_Update/ack
      -- 
    ack_7584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2886_delayed_1_0_3000_inst_ack_1, ack => convolve_CP_6623_elements(297)); -- 
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	224 
    -- CP-element group 298: 	228 
    -- CP-element group 298: 	232 
    -- CP-element group 298: 	236 
    -- CP-element group 298: 	220 
    -- CP-element group 298: 	160 
    -- CP-element group 298: 	164 
    -- CP-element group 298: 	168 
    -- CP-element group 298: 	172 
    -- CP-element group 298: 	156 
    -- CP-element group 298: 	180 
    -- CP-element group 298: 	184 
    -- CP-element group 298: 	188 
    -- CP-element group 298: 	256 
    -- CP-element group 298: 	260 
    -- CP-element group 298: 	144 
    -- CP-element group 298: 	148 
    -- CP-element group 298: 	152 
    -- CP-element group 298: 	240 
    -- CP-element group 298: 	244 
    -- CP-element group 298: 	248 
    -- CP-element group 298: 	252 
    -- CP-element group 298: 	176 
    -- CP-element group 298: 	297 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_Sample/rr
      -- 
    rr_7592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(298), ack => CONCAT_u8_u16_3009_inst_req_0); -- 
    convolve_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 24) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1);
      constant place_markings: IntegerArray(0 to 24)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 1);
      constant place_delays: IntegerArray(0 to 24) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 25); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(224) & convolve_CP_6623_elements(228) & convolve_CP_6623_elements(232) & convolve_CP_6623_elements(236) & convolve_CP_6623_elements(220) & convolve_CP_6623_elements(160) & convolve_CP_6623_elements(164) & convolve_CP_6623_elements(168) & convolve_CP_6623_elements(172) & convolve_CP_6623_elements(156) & convolve_CP_6623_elements(180) & convolve_CP_6623_elements(184) & convolve_CP_6623_elements(188) & convolve_CP_6623_elements(256) & convolve_CP_6623_elements(260) & convolve_CP_6623_elements(144) & convolve_CP_6623_elements(148) & convolve_CP_6623_elements(152) & convolve_CP_6623_elements(240) & convolve_CP_6623_elements(244) & convolve_CP_6623_elements(248) & convolve_CP_6623_elements(252) & convolve_CP_6623_elements(176) & convolve_CP_6623_elements(297) & convolve_CP_6623_elements(300);
      gj_convolve_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 25, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: marked-predecessors 
    -- CP-element group 299: 	301 
    -- CP-element group 299: 	303 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	301 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_update_start_
      -- CP-element group 299: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_Update/cr
      -- 
    cr_7597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(299), ack => CONCAT_u8_u16_3009_inst_req_1); -- 
    convolve_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(301) & convolve_CP_6623_elements(303);
      gj_convolve_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	226 
    -- CP-element group 300: 	230 
    -- CP-element group 300: 	234 
    -- CP-element group 300: 	238 
    -- CP-element group 300: 	218 
    -- CP-element group 300: 	222 
    -- CP-element group 300: 	162 
    -- CP-element group 300: 	166 
    -- CP-element group 300: 	170 
    -- CP-element group 300: 	154 
    -- CP-element group 300: 	158 
    -- CP-element group 300: 	182 
    -- CP-element group 300: 	186 
    -- CP-element group 300: 	254 
    -- CP-element group 300: 	258 
    -- CP-element group 300: 	142 
    -- CP-element group 300: 	146 
    -- CP-element group 300: 	150 
    -- CP-element group 300: 	242 
    -- CP-element group 300: 	246 
    -- CP-element group 300: 	250 
    -- CP-element group 300: 	174 
    -- CP-element group 300: 	178 
    -- CP-element group 300: 	295 
    -- CP-element group 300: 	298 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_Sample/ra
      -- 
    ra_7593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_3009_inst_ack_0, ack => convolve_CP_6623_elements(300)); -- 
    -- CP-element group 301:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	299 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301: marked-successors 
    -- CP-element group 301: 	299 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/CONCAT_u8_u16_3009_Update/ca
      -- 
    ca_7598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_3009_inst_ack_1, ack => convolve_CP_6623_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	297 
    -- CP-element group 302: 	301 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	304 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_Sample/req
      -- 
    req_7606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(302), ack => WPIPE_output_pipe_3004_inst_req_0); -- 
    convolve_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(297) & convolve_CP_6623_elements(301) & convolve_CP_6623_elements(304);
      gj_convolve_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	295 
    -- CP-element group 303: 	299 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_update_start_
      -- CP-element group 303: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_Update/req
      -- 
    ack_7607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3004_inst_ack_0, ack => convolve_CP_6623_elements(303)); -- 
    req_7611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(303), ack => WPIPE_output_pipe_3004_inst_req_1); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	306 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	302 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/WPIPE_output_pipe_3004_Update/ack
      -- 
    ack_7612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3004_inst_ack_1, ack => convolve_CP_6623_elements(304)); -- 
    -- CP-element group 305:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	23 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	24 
    -- CP-element group 305:  members (1) 
      -- CP-element group 305: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_6623_elements(305) is a control-delay.
    cp_element_305_delay: control_delay_element  generic map(name => " 305_delay", delay_value => 1)  port map(req => convolve_CP_6623_elements(23), ack => convolve_CP_6623_elements(305), clk => clk, reset =>reset);
    -- CP-element group 306:  join  transition  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	195 
    -- CP-element group 306: 	216 
    -- CP-element group 306: 	26 
    -- CP-element group 306: 	202 
    -- CP-element group 306: 	209 
    -- CP-element group 306: 	271 
    -- CP-element group 306: 	278 
    -- CP-element group 306: 	285 
    -- CP-element group 306: 	289 
    -- CP-element group 306: 	293 
    -- CP-element group 306: 	304 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	20 
    -- CP-element group 306:  members (1) 
      -- CP-element group 306: 	 branch_block_stmt_2566/do_while_stmt_2583/do_while_stmt_2583_loop_body/$exit
      -- 
    convolve_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolve_CP_6623_elements(195) & convolve_CP_6623_elements(216) & convolve_CP_6623_elements(26) & convolve_CP_6623_elements(202) & convolve_CP_6623_elements(209) & convolve_CP_6623_elements(271) & convolve_CP_6623_elements(278) & convolve_CP_6623_elements(285) & convolve_CP_6623_elements(289) & convolve_CP_6623_elements(293) & convolve_CP_6623_elements(304);
      gj_convolve_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6623_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	19 
    -- CP-element group 307: successors 
    -- CP-element group 307:  members (2) 
      -- CP-element group 307: 	 branch_block_stmt_2566/do_while_stmt_2583/loop_exit/$exit
      -- CP-element group 307: 	 branch_block_stmt_2566/do_while_stmt_2583/loop_exit/ack
      -- 
    ack_7617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2583_branch_ack_0, ack => convolve_CP_6623_elements(307)); -- 
    -- CP-element group 308:  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	19 
    -- CP-element group 308: successors 
    -- CP-element group 308:  members (2) 
      -- CP-element group 308: 	 branch_block_stmt_2566/do_while_stmt_2583/loop_taken/$exit
      -- CP-element group 308: 	 branch_block_stmt_2566/do_while_stmt_2583/loop_taken/ack
      -- 
    ack_7621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2583_branch_ack_1, ack => convolve_CP_6623_elements(308)); -- 
    -- CP-element group 309:  transition  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	17 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	2 
    -- CP-element group 309:  members (1) 
      -- CP-element group 309: 	 branch_block_stmt_2566/do_while_stmt_2583/$exit
      -- 
    convolve_CP_6623_elements(309) <= convolve_CP_6623_elements(17);
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	2 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_update_start_
      -- CP-element group 310: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_Sample/ack
      -- CP-element group 310: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_Update/req
      -- 
    ack_7634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3014_inst_ack_0, ack => convolve_CP_6623_elements(310)); -- 
    req_7638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(310), ack => WPIPE_input_done_pipe_3014_inst_req_1); -- 
    -- CP-element group 311:  transition  place  input  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (8) 
      -- CP-element group 311: 	 branch_block_stmt_2566/loopback
      -- CP-element group 311: 	 branch_block_stmt_2566/assign_stmt_3016__exit__
      -- CP-element group 311: 	 branch_block_stmt_2566/assign_stmt_3016/$exit
      -- CP-element group 311: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_2566/assign_stmt_3016/WPIPE_input_done_pipe_3014_Update/ack
      -- CP-element group 311: 	 branch_block_stmt_2566/loopback_PhiReq/$entry
      -- CP-element group 311: 	 branch_block_stmt_2566/loopback_PhiReq/$exit
      -- 
    ack_7639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3014_inst_ack_1, ack => convolve_CP_6623_elements(311)); -- 
    -- CP-element group 312:  merge  fork  transition  place  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	0 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	3 
    -- CP-element group 312: 	14 
    -- CP-element group 312: 	10 
    -- CP-element group 312: 	11 
    -- CP-element group 312: 	6 
    -- CP-element group 312:  members (22) 
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582__entry__
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_2566/merge_stmt_2567__exit__
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_update_start_
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_update_start_
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_Sample/rr
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2576_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_Update/cr
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2581_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/$entry
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_size_pipe_2579_Sample/rr
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/SUB_u16_u16_2571_update_start_
      -- CP-element group 312: 	 branch_block_stmt_2566/assign_stmt_2572_to_assign_stmt_2582/RPIPE_num_out_pipe_2569_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_2566/merge_stmt_2567_PhiReqMerge
      -- CP-element group 312: 	 branch_block_stmt_2566/merge_stmt_2567_PhiAck/$entry
      -- CP-element group 312: 	 branch_block_stmt_2566/merge_stmt_2567_PhiAck/$exit
      -- CP-element group 312: 	 branch_block_stmt_2566/merge_stmt_2567_PhiAck/dummy
      -- 
    cr_6725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(312), ack => SUB_u16_u16_2581_inst_req_1); -- 
    cr_6697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(312), ack => SUB_u16_u16_2576_inst_req_1); -- 
    rr_6654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(312), ack => RPIPE_num_out_pipe_2569_inst_req_0); -- 
    cr_6669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(312), ack => SUB_u16_u16_2571_inst_req_1); -- 
    rr_6710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6623_elements(312), ack => RPIPE_size_pipe_2579_inst_req_0); -- 
    convolve_CP_6623_elements(312) <= OrReduce(convolve_CP_6623_elements(0) & convolve_CP_6623_elements(311));
    convolve_do_while_stmt_2583_terminator_7622: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_2583_terminator_7622", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_6623_elements(20),loop_continue => convolve_CP_6623_elements(308),loop_terminate => convolve_CP_6623_elements(307),loop_back => convolve_CP_6623_elements(18),loop_exit => convolve_CP_6623_elements(17),clk => clk, reset => reset); -- 
    phi_stmt_2585_phi_seq_6790_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6623_elements(35);
      convolve_CP_6623_elements(38)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6623_elements(38);
      convolve_CP_6623_elements(39)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6623_elements(40);
      convolve_CP_6623_elements(36) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6623_elements(33);
      convolve_CP_6623_elements(42)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6623_elements(44);
      convolve_CP_6623_elements(43)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6623_elements(45);
      convolve_CP_6623_elements(34) <= phi_mux_reqs(1);
      phi_stmt_2585_phi_seq_6790 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2585_phi_seq_6790") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6623_elements(25), 
          phi_sample_ack => convolve_CP_6623_elements(31), 
          phi_update_req => convolve_CP_6623_elements(27), 
          phi_update_ack => convolve_CP_6623_elements(32), 
          phi_mux_ack => convolve_CP_6623_elements(37), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2591_phi_seq_6834_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6623_elements(54);
      convolve_CP_6623_elements(57)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6623_elements(57);
      convolve_CP_6623_elements(58)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6623_elements(59);
      convolve_CP_6623_elements(55) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6623_elements(52);
      convolve_CP_6623_elements(61)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6623_elements(63);
      convolve_CP_6623_elements(62)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6623_elements(64);
      convolve_CP_6623_elements(53) <= phi_mux_reqs(1);
      phi_stmt_2591_phi_seq_6834 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2591_phi_seq_6834") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6623_elements(48), 
          phi_sample_ack => convolve_CP_6623_elements(49), 
          phi_update_req => convolve_CP_6623_elements(50), 
          phi_update_ack => convolve_CP_6623_elements(51), 
          phi_mux_ack => convolve_CP_6623_elements(56), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2596_phi_seq_6878_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6623_elements(73);
      convolve_CP_6623_elements(76)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6623_elements(76);
      convolve_CP_6623_elements(77)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6623_elements(78);
      convolve_CP_6623_elements(74) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6623_elements(71);
      convolve_CP_6623_elements(80)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6623_elements(82);
      convolve_CP_6623_elements(81)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6623_elements(83);
      convolve_CP_6623_elements(72) <= phi_mux_reqs(1);
      phi_stmt_2596_phi_seq_6878 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2596_phi_seq_6878") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6623_elements(67), 
          phi_sample_ack => convolve_CP_6623_elements(68), 
          phi_update_req => convolve_CP_6623_elements(69), 
          phi_update_ack => convolve_CP_6623_elements(70), 
          phi_mux_ack => convolve_CP_6623_elements(75), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2601_phi_seq_6922_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6623_elements(92);
      convolve_CP_6623_elements(95)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6623_elements(95);
      convolve_CP_6623_elements(96)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6623_elements(97);
      convolve_CP_6623_elements(93) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6623_elements(90);
      convolve_CP_6623_elements(99)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6623_elements(101);
      convolve_CP_6623_elements(100)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6623_elements(102);
      convolve_CP_6623_elements(91) <= phi_mux_reqs(1);
      phi_stmt_2601_phi_seq_6922 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2601_phi_seq_6922") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6623_elements(86), 
          phi_sample_ack => convolve_CP_6623_elements(87), 
          phi_update_req => convolve_CP_6623_elements(88), 
          phi_update_ack => convolve_CP_6623_elements(89), 
          phi_mux_ack => convolve_CP_6623_elements(94), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2606_phi_seq_6966_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6623_elements(111);
      convolve_CP_6623_elements(114)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6623_elements(114);
      convolve_CP_6623_elements(115)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6623_elements(116);
      convolve_CP_6623_elements(112) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6623_elements(109);
      convolve_CP_6623_elements(118)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6623_elements(120);
      convolve_CP_6623_elements(119)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6623_elements(121);
      convolve_CP_6623_elements(110) <= phi_mux_reqs(1);
      phi_stmt_2606_phi_seq_6966 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2606_phi_seq_6966") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6623_elements(105), 
          phi_sample_ack => convolve_CP_6623_elements(106), 
          phi_update_req => convolve_CP_6623_elements(107), 
          phi_update_ack => convolve_CP_6623_elements(108), 
          phi_mux_ack => convolve_CP_6623_elements(113), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2612_phi_seq_7010_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6623_elements(130);
      convolve_CP_6623_elements(133)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6623_elements(133);
      convolve_CP_6623_elements(134)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6623_elements(135);
      convolve_CP_6623_elements(131) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6623_elements(128);
      convolve_CP_6623_elements(137)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6623_elements(139);
      convolve_CP_6623_elements(138)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6623_elements(140);
      convolve_CP_6623_elements(129) <= phi_mux_reqs(1);
      phi_stmt_2612_phi_seq_7010 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2612_phi_seq_7010") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6623_elements(124), 
          phi_sample_ack => convolve_CP_6623_elements(125), 
          phi_update_req => convolve_CP_6623_elements(126), 
          phi_update_ack => convolve_CP_6623_elements(127), 
          phi_mux_ack => convolve_CP_6623_elements(132), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_6742_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_6623_elements(21);
        preds(1)  <= convolve_CP_6623_elements(22);
        entry_tmerge_6742 : transition_merge -- 
          generic map(name => " entry_tmerge_6742")
          port map (preds => preds, symbol_out => convolve_CP_6623_elements(23));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_i8_i8_2862_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2865_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2874_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2877_wire : std_logic_vector(7 downto 0);
    signal ADD_u16_u16_2949_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2969_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2978_wire : std_logic_vector(15 downto 0);
    signal ADD_u2_u2_2958_wire : std_logic_vector(1 downto 0);
    signal AND_u1_u1_2915_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u8_u16_3009_wire : std_logic_vector(15 downto 0);
    signal EQ_u16_u1_2621_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2751_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2754_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2624_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2888_wire : std_logic_vector(0 downto 0);
    signal MUL_i8_i8_2823_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2829_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2835_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2841_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2847_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2853_wire : std_logic_vector(7 downto 0);
    signal MUX_2959_wire : std_logic_vector(1 downto 0);
    signal MUX_2970_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_3013_wire : std_logic_vector(0 downto 0);
    signal RPIPE_num_out_pipe_2569_wire : std_logic_vector(15 downto 0);
    signal RPIPE_num_out_pipe_2574_wire : std_logic_vector(15 downto 0);
    signal RPIPE_size_pipe_2579_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_2810_2810_delayed_1_0_2906 : std_logic_vector(15 downto 0);
    signal UGT_u2_u1_2701_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_2698_wire : std_logic_vector(0 downto 0);
    signal acc1_2585 : std_logic_vector(7 downto 0);
    signal acc1_2767_delayed_1_0_2858 : std_logic_vector(7 downto 0);
    signal acc2_2591 : std_logic_vector(7 downto 0);
    signal acc2_2776_delayed_1_0_2870 : std_logic_vector(7 downto 0);
    signal acc_val1_2867 : std_logic_vector(7 downto 0);
    signal acc_val2_2879 : std_logic_vector(7 downto 0);
    signal all_done_flag_2922 : std_logic_vector(0 downto 0);
    signal chl_2612 : std_logic_vector(15 downto 0);
    signal chl_done_2884 : std_logic_vector(0 downto 0);
    signal col_2601 : std_logic_vector(15 downto 0);
    signal col_done_2896 : std_logic_vector(0 downto 0);
    signal iread1_2667 : std_logic_vector(7 downto 0);
    signal iread2_2676 : std_logic_vector(7 downto 0);
    signal iread3_2685 : std_logic_vector(7 downto 0);
    signal iread4_2694 : std_logic_vector(7 downto 0);
    signal ival1_2735 : std_logic_vector(7 downto 0);
    signal ival2_2739 : std_logic_vector(7 downto 0);
    signal ival3_2743 : std_logic_vector(7 downto 0);
    signal ival4_2747 : std_logic_vector(7 downto 0);
    signal konst_2570_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2575_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2580_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2620_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2623_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2700_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2750_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2753_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2887_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2904_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2946_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2948_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2955_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2957_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2966_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2968_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2977_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2987_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2996_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3015_wire_constant : std_logic_vector(7 downto 0);
    signal kread1_2789 : std_logic_vector(7 downto 0);
    signal kread2_2798 : std_logic_vector(7 downto 0);
    signal kread3_2807 : std_logic_vector(7 downto 0);
    signal kval1_2811 : std_logic_vector(7 downto 0);
    signal kval2_2815 : std_logic_vector(7 downto 0);
    signal kval3_2819 : std_logic_vector(7 downto 0);
    signal mul_val1_2825 : std_logic_vector(7 downto 0);
    signal mul_val2_2831 : std_logic_vector(7 downto 0);
    signal mul_val3_2837 : std_logic_vector(7 downto 0);
    signal mul_val4_2843 : std_logic_vector(7 downto 0);
    signal mul_val5_2849 : std_logic_vector(7 downto 0);
    signal mul_val6_2855 : std_logic_vector(7 downto 0);
    signal n_chl_2951 : std_logic_vector(15 downto 0);
    signal n_chl_2951_2616_buffered : std_logic_vector(15 downto 0);
    signal n_col_2973 : std_logic_vector(15 downto 0);
    signal n_col_2973_2605_buffered : std_logic_vector(15 downto 0);
    signal n_num_2962 : std_logic_vector(1 downto 0);
    signal n_num_2962_2611_buffered : std_logic_vector(1 downto 0);
    signal n_row_2981 : std_logic_vector(15 downto 0);
    signal n_row_2981_2600_buffered : std_logic_vector(15 downto 0);
    signal nacc1_2990 : std_logic_vector(7 downto 0);
    signal nacc1_2990_2590_buffered : std_logic_vector(7 downto 0);
    signal nacc2_2999 : std_logic_vector(7 downto 0);
    signal nacc2_2999_2595_buffered : std_logic_vector(7 downto 0);
    signal num_2606 : std_logic_vector(1 downto 0);
    signal num_chl_2582 : std_logic_vector(15 downto 0);
    signal num_col_2577 : std_logic_vector(15 downto 0);
    signal num_done_2875_delayed_1_0_2984 : std_logic_vector(0 downto 0);
    signal num_done_2881_delayed_1_0_2993 : std_logic_vector(0 downto 0);
    signal num_done_2886_delayed_1_0_3002 : std_logic_vector(0 downto 0);
    signal num_done_2891 : std_logic_vector(0 downto 0);
    signal num_row_2572 : std_logic_vector(15 downto 0);
    signal out_done_flag_2911 : std_logic_vector(0 downto 0);
    signal read_ip_2603_delayed_1_0_2661 : std_logic_vector(0 downto 0);
    signal read_ip_2609_delayed_1_0_2670 : std_logic_vector(0 downto 0);
    signal read_ip_2615_delayed_1_0_2679 : std_logic_vector(0 downto 0);
    signal read_ip_2621_delayed_1_0_2688 : std_logic_vector(0 downto 0);
    signal read_ip_2626 : std_logic_vector(0 downto 0);
    signal read_k_2701_delayed_1_0_2783 : std_logic_vector(0 downto 0);
    signal read_k_2707_delayed_1_0_2792 : std_logic_vector(0 downto 0);
    signal read_k_2713_delayed_1_0_2801 : std_logic_vector(0 downto 0);
    signal read_k_2756 : std_logic_vector(0 downto 0);
    signal row_2596 : std_logic_vector(15 downto 0);
    signal row_done_2901 : std_logic_vector(0 downto 0);
    signal store_kernel_2824_delayed_1_0_2925 : std_logic_vector(0 downto 0);
    signal store_kernel_2828_delayed_1_0_2932 : std_logic_vector(0 downto 0);
    signal store_kernel_2832_delayed_1_0_2939 : std_logic_vector(0 downto 0);
    signal store_kernel_2917 : std_logic_vector(0 downto 0);
    signal temp1_1_2646 : std_logic_vector(7 downto 0);
    signal temp1_2_2650 : std_logic_vector(7 downto 0);
    signal temp1_3_2654 : std_logic_vector(7 downto 0);
    signal temp1_4_2658 : std_logic_vector(7 downto 0);
    signal temp2_1_2630 : std_logic_vector(7 downto 0);
    signal temp2_2_2634 : std_logic_vector(7 downto 0);
    signal temp2_3_2638 : std_logic_vector(7 downto 0);
    signal temp2_4_2642 : std_logic_vector(7 downto 0);
    signal tempk1_1_2760 : std_logic_vector(7 downto 0);
    signal tempk1_2_2764 : std_logic_vector(7 downto 0);
    signal tempk1_3_2768 : std_logic_vector(7 downto 0);
    signal tempk2_1_2772 : std_logic_vector(7 downto 0);
    signal tempk2_2_2776 : std_logic_vector(7 downto 0);
    signal tempk2_3_2780 : std_logic_vector(7 downto 0);
    signal type_cast_2589_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2594_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2599_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2604_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2610_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_2615_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3006_wire : std_logic_vector(7 downto 0);
    signal type_cast_3008_wire : std_logic_vector(7 downto 0);
    signal write_input_2635_delayed_1_0_2706 : std_logic_vector(0 downto 0);
    signal write_input_2639_delayed_1_0_2713 : std_logic_vector(0 downto 0);
    signal write_input_2643_delayed_1_0_2720 : std_logic_vector(0 downto 0);
    signal write_input_2647_delayed_1_0_2727 : std_logic_vector(0 downto 0);
    signal write_input_2703 : std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip4
    signal xxconvolvexxconv_ip4_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_ip4_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip4_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip4
    signal xxconvolvexxconv_ip4_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_ip4_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip4_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_2570_wire_constant <= "0000000000000001";
    konst_2575_wire_constant <= "0000000000000001";
    konst_2580_wire_constant <= "0000000000000001";
    konst_2620_wire_constant <= "0000000000000000";
    konst_2623_wire_constant <= "10";
    konst_2700_wire_constant <= "00";
    konst_2750_wire_constant <= "0000000000000000";
    konst_2753_wire_constant <= "0000000000000000";
    konst_2887_wire_constant <= "10";
    konst_2904_wire_constant <= "0000000000000001";
    konst_2946_wire_constant <= "0000000000000000";
    konst_2948_wire_constant <= "0000000000000001";
    konst_2955_wire_constant <= "00";
    konst_2957_wire_constant <= "01";
    konst_2966_wire_constant <= "0000000000000000";
    konst_2968_wire_constant <= "0000000000000001";
    konst_2977_wire_constant <= "0000000000000010";
    konst_2987_wire_constant <= "00000000";
    konst_2996_wire_constant <= "00000000";
    konst_3015_wire_constant <= "00000001";
    type_cast_2589_wire_constant <= "00000000";
    type_cast_2594_wire_constant <= "00000000";
    type_cast_2599_wire_constant <= "0000000000000000";
    type_cast_2604_wire_constant <= "0000000000000000";
    type_cast_2610_wire_constant <= "00";
    type_cast_2615_wire_constant <= "0000000000000000";
    phi_stmt_2585: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2589_wire_constant & nacc1_2990_2590_buffered;
      req <= phi_stmt_2585_req_0 & phi_stmt_2585_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2585",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2585_ack_0,
          idata => idata,
          odata => acc1_2585,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2585
    phi_stmt_2591: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2594_wire_constant & nacc2_2999_2595_buffered;
      req <= phi_stmt_2591_req_0 & phi_stmt_2591_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2591",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2591_ack_0,
          idata => idata,
          odata => acc2_2591,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2591
    phi_stmt_2596: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2599_wire_constant & n_row_2981_2600_buffered;
      req <= phi_stmt_2596_req_0 & phi_stmt_2596_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2596",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2596_ack_0,
          idata => idata,
          odata => row_2596,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2596
    phi_stmt_2601: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2604_wire_constant & n_col_2973_2605_buffered;
      req <= phi_stmt_2601_req_0 & phi_stmt_2601_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2601",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2601_ack_0,
          idata => idata,
          odata => col_2601,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2601
    phi_stmt_2606: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2610_wire_constant & n_num_2962_2611_buffered;
      req <= phi_stmt_2606_req_0 & phi_stmt_2606_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2606",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2606_ack_0,
          idata => idata,
          odata => num_2606,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2606
    phi_stmt_2612: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2615_wire_constant & n_chl_2951_2616_buffered;
      req <= phi_stmt_2612_req_0 & phi_stmt_2612_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2612",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2612_ack_0,
          idata => idata,
          odata => chl_2612,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2612
    -- flow-through select operator MUX_2666_inst
    iread1_2667 <= temp2_1_2630 when (read_ip_2603_delayed_1_0_2661(0) /=  '0') else temp1_1_2646;
    -- flow-through select operator MUX_2675_inst
    iread2_2676 <= temp2_2_2634 when (read_ip_2609_delayed_1_0_2670(0) /=  '0') else temp1_2_2650;
    -- flow-through select operator MUX_2684_inst
    iread3_2685 <= temp2_3_2638 when (read_ip_2615_delayed_1_0_2679(0) /=  '0') else temp1_3_2654;
    -- flow-through select operator MUX_2693_inst
    iread4_2694 <= temp2_4_2642 when (read_ip_2621_delayed_1_0_2688(0) /=  '0') else temp1_4_2658;
    -- flow-through select operator MUX_2788_inst
    kread1_2789 <= tempk1_1_2760 when (read_k_2701_delayed_1_0_2783(0) /=  '0') else tempk2_1_2772;
    -- flow-through select operator MUX_2797_inst
    kread2_2798 <= tempk1_2_2764 when (read_k_2707_delayed_1_0_2792(0) /=  '0') else tempk2_2_2776;
    -- flow-through select operator MUX_2806_inst
    kread3_2807 <= tempk1_3_2768 when (read_k_2713_delayed_1_0_2801(0) /=  '0') else tempk2_3_2780;
    -- flow-through select operator MUX_2950_inst
    n_chl_2951 <= konst_2946_wire_constant when (chl_done_2884(0) /=  '0') else ADD_u16_u16_2949_wire;
    -- flow-through select operator MUX_2959_inst
    MUX_2959_wire <= konst_2955_wire_constant when (num_done_2891(0) /=  '0') else ADD_u2_u2_2958_wire;
    -- flow-through select operator MUX_2961_inst
    n_num_2962 <= MUX_2959_wire when (chl_done_2884(0) /=  '0') else num_2606;
    -- flow-through select operator MUX_2970_inst
    MUX_2970_wire <= konst_2966_wire_constant when (col_done_2896(0) /=  '0') else ADD_u16_u16_2969_wire;
    -- flow-through select operator MUX_2972_inst
    n_col_2973 <= MUX_2970_wire when (num_done_2891(0) /=  '0') else col_2601;
    -- flow-through select operator MUX_2980_inst
    n_row_2981 <= ADD_u16_u16_2978_wire when (row_done_2901(0) /=  '0') else row_2596;
    -- flow-through select operator MUX_2989_inst
    nacc1_2990 <= konst_2987_wire_constant when (num_done_2875_delayed_1_0_2984(0) /=  '0') else acc_val1_2867;
    -- flow-through select operator MUX_2998_inst
    nacc2_2999 <= konst_2996_wire_constant when (num_done_2881_delayed_1_0_2993(0) /=  '0') else acc_val2_2879;
    W_acc1_2767_delayed_1_0_2856_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc1_2767_delayed_1_0_2856_inst_req_0;
      W_acc1_2767_delayed_1_0_2856_inst_ack_0<= wack(0);
      rreq(0) <= W_acc1_2767_delayed_1_0_2856_inst_req_1;
      W_acc1_2767_delayed_1_0_2856_inst_ack_1<= rack(0);
      W_acc1_2767_delayed_1_0_2856_inst : InterlockBuffer generic map ( -- 
        name => "W_acc1_2767_delayed_1_0_2856_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc1_2585,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc1_2767_delayed_1_0_2858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_acc2_2776_delayed_1_0_2868_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc2_2776_delayed_1_0_2868_inst_req_0;
      W_acc2_2776_delayed_1_0_2868_inst_ack_0<= wack(0);
      rreq(0) <= W_acc2_2776_delayed_1_0_2868_inst_req_1;
      W_acc2_2776_delayed_1_0_2868_inst_ack_1<= rack(0);
      W_acc2_2776_delayed_1_0_2868_inst : InterlockBuffer generic map ( -- 
        name => "W_acc2_2776_delayed_1_0_2868_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc2_2591,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc2_2776_delayed_1_0_2870,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2875_delayed_1_0_2982_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2875_delayed_1_0_2982_inst_req_0;
      W_num_done_2875_delayed_1_0_2982_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2875_delayed_1_0_2982_inst_req_1;
      W_num_done_2875_delayed_1_0_2982_inst_ack_1<= rack(0);
      W_num_done_2875_delayed_1_0_2982_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2875_delayed_1_0_2982_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2891,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2875_delayed_1_0_2984,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2881_delayed_1_0_2991_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2881_delayed_1_0_2991_inst_req_0;
      W_num_done_2881_delayed_1_0_2991_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2881_delayed_1_0_2991_inst_req_1;
      W_num_done_2881_delayed_1_0_2991_inst_ack_1<= rack(0);
      W_num_done_2881_delayed_1_0_2991_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2881_delayed_1_0_2991_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2891,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2881_delayed_1_0_2993,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2886_delayed_1_0_3000_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2886_delayed_1_0_3000_inst_req_0;
      W_num_done_2886_delayed_1_0_3000_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2886_delayed_1_0_3000_inst_req_1;
      W_num_done_2886_delayed_1_0_3000_inst_ack_1<= rack(0);
      W_num_done_2886_delayed_1_0_3000_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2886_delayed_1_0_3000_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2891,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2886_delayed_1_0_3002,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2603_delayed_1_0_2659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2603_delayed_1_0_2659_inst_req_0;
      W_read_ip_2603_delayed_1_0_2659_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2603_delayed_1_0_2659_inst_req_1;
      W_read_ip_2603_delayed_1_0_2659_inst_ack_1<= rack(0);
      W_read_ip_2603_delayed_1_0_2659_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2603_delayed_1_0_2659_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2603_delayed_1_0_2661,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2609_delayed_1_0_2668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2609_delayed_1_0_2668_inst_req_0;
      W_read_ip_2609_delayed_1_0_2668_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2609_delayed_1_0_2668_inst_req_1;
      W_read_ip_2609_delayed_1_0_2668_inst_ack_1<= rack(0);
      W_read_ip_2609_delayed_1_0_2668_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2609_delayed_1_0_2668_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2609_delayed_1_0_2670,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2615_delayed_1_0_2677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2615_delayed_1_0_2677_inst_req_0;
      W_read_ip_2615_delayed_1_0_2677_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2615_delayed_1_0_2677_inst_req_1;
      W_read_ip_2615_delayed_1_0_2677_inst_ack_1<= rack(0);
      W_read_ip_2615_delayed_1_0_2677_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2615_delayed_1_0_2677_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2615_delayed_1_0_2679,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2621_delayed_1_0_2686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2621_delayed_1_0_2686_inst_req_0;
      W_read_ip_2621_delayed_1_0_2686_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2621_delayed_1_0_2686_inst_req_1;
      W_read_ip_2621_delayed_1_0_2686_inst_ack_1<= rack(0);
      W_read_ip_2621_delayed_1_0_2686_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2621_delayed_1_0_2686_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2621_delayed_1_0_2688,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2701_delayed_1_0_2781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2701_delayed_1_0_2781_inst_req_0;
      W_read_k_2701_delayed_1_0_2781_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2701_delayed_1_0_2781_inst_req_1;
      W_read_k_2701_delayed_1_0_2781_inst_ack_1<= rack(0);
      W_read_k_2701_delayed_1_0_2781_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2701_delayed_1_0_2781_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2701_delayed_1_0_2783,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2707_delayed_1_0_2790_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2707_delayed_1_0_2790_inst_req_0;
      W_read_k_2707_delayed_1_0_2790_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2707_delayed_1_0_2790_inst_req_1;
      W_read_k_2707_delayed_1_0_2790_inst_ack_1<= rack(0);
      W_read_k_2707_delayed_1_0_2790_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2707_delayed_1_0_2790_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2707_delayed_1_0_2792,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2713_delayed_1_0_2799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2713_delayed_1_0_2799_inst_req_0;
      W_read_k_2713_delayed_1_0_2799_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2713_delayed_1_0_2799_inst_req_1;
      W_read_k_2713_delayed_1_0_2799_inst_ack_1<= rack(0);
      W_read_k_2713_delayed_1_0_2799_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2713_delayed_1_0_2799_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2713_delayed_1_0_2801,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2824_delayed_1_0_2923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2824_delayed_1_0_2923_inst_req_0;
      W_store_kernel_2824_delayed_1_0_2923_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2824_delayed_1_0_2923_inst_req_1;
      W_store_kernel_2824_delayed_1_0_2923_inst_ack_1<= rack(0);
      W_store_kernel_2824_delayed_1_0_2923_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2824_delayed_1_0_2923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2824_delayed_1_0_2925,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2828_delayed_1_0_2930_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2828_delayed_1_0_2930_inst_req_0;
      W_store_kernel_2828_delayed_1_0_2930_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2828_delayed_1_0_2930_inst_req_1;
      W_store_kernel_2828_delayed_1_0_2930_inst_ack_1<= rack(0);
      W_store_kernel_2828_delayed_1_0_2930_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2828_delayed_1_0_2930_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2828_delayed_1_0_2932,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2832_delayed_1_0_2937_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2832_delayed_1_0_2937_inst_req_0;
      W_store_kernel_2832_delayed_1_0_2937_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2832_delayed_1_0_2937_inst_req_1;
      W_store_kernel_2832_delayed_1_0_2937_inst_ack_1<= rack(0);
      W_store_kernel_2832_delayed_1_0_2937_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2832_delayed_1_0_2937_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2832_delayed_1_0_2939,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2635_delayed_1_0_2704_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2635_delayed_1_0_2704_inst_req_0;
      W_write_input_2635_delayed_1_0_2704_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2635_delayed_1_0_2704_inst_req_1;
      W_write_input_2635_delayed_1_0_2704_inst_ack_1<= rack(0);
      W_write_input_2635_delayed_1_0_2704_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2635_delayed_1_0_2704_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2635_delayed_1_0_2706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2639_delayed_1_0_2711_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2639_delayed_1_0_2711_inst_req_0;
      W_write_input_2639_delayed_1_0_2711_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2639_delayed_1_0_2711_inst_req_1;
      W_write_input_2639_delayed_1_0_2711_inst_ack_1<= rack(0);
      W_write_input_2639_delayed_1_0_2711_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2639_delayed_1_0_2711_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2639_delayed_1_0_2713,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2643_delayed_1_0_2718_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2643_delayed_1_0_2718_inst_req_0;
      W_write_input_2643_delayed_1_0_2718_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2643_delayed_1_0_2718_inst_req_1;
      W_write_input_2643_delayed_1_0_2718_inst_ack_1<= rack(0);
      W_write_input_2643_delayed_1_0_2718_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2643_delayed_1_0_2718_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2643_delayed_1_0_2720,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2647_delayed_1_0_2725_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2647_delayed_1_0_2725_inst_req_0;
      W_write_input_2647_delayed_1_0_2725_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2647_delayed_1_0_2725_inst_req_1;
      W_write_input_2647_delayed_1_0_2725_inst_ack_1<= rack(0);
      W_write_input_2647_delayed_1_0_2725_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2647_delayed_1_0_2725_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2647_delayed_1_0_2727,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_2951_2616_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_2951_2616_buf_req_0;
      n_chl_2951_2616_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_2951_2616_buf_req_1;
      n_chl_2951_2616_buf_ack_1<= rack(0);
      n_chl_2951_2616_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_2951_2616_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_2951,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_2951_2616_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_2973_2605_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_2973_2605_buf_req_0;
      n_col_2973_2605_buf_ack_0<= wack(0);
      rreq(0) <= n_col_2973_2605_buf_req_1;
      n_col_2973_2605_buf_ack_1<= rack(0);
      n_col_2973_2605_buf : InterlockBuffer generic map ( -- 
        name => "n_col_2973_2605_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_2973,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_2973_2605_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_num_2962_2611_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_num_2962_2611_buf_req_0;
      n_num_2962_2611_buf_ack_0<= wack(0);
      rreq(0) <= n_num_2962_2611_buf_req_1;
      n_num_2962_2611_buf_ack_1<= rack(0);
      n_num_2962_2611_buf : InterlockBuffer generic map ( -- 
        name => "n_num_2962_2611_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_num_2962,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_num_2962_2611_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_2981_2600_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_2981_2600_buf_req_0;
      n_row_2981_2600_buf_ack_0<= wack(0);
      rreq(0) <= n_row_2981_2600_buf_req_1;
      n_row_2981_2600_buf_ack_1<= rack(0);
      n_row_2981_2600_buf : InterlockBuffer generic map ( -- 
        name => "n_row_2981_2600_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_2981,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_2981_2600_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc1_2990_2590_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc1_2990_2590_buf_req_0;
      nacc1_2990_2590_buf_ack_0<= wack(0);
      rreq(0) <= nacc1_2990_2590_buf_req_1;
      nacc1_2990_2590_buf_ack_1<= rack(0);
      nacc1_2990_2590_buf : InterlockBuffer generic map ( -- 
        name => "nacc1_2990_2590_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc1_2990,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc1_2990_2590_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc2_2999_2595_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc2_2999_2595_buf_req_0;
      nacc2_2999_2595_buf_ack_0<= wack(0);
      rreq(0) <= nacc2_2999_2595_buf_req_1;
      nacc2_2999_2595_buf_ack_1<= rack(0);
      nacc2_2999_2595_buf : InterlockBuffer generic map ( -- 
        name => "nacc2_2999_2595_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc2_2999,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc2_2999_2595_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2734_inst
    process(iread1_2667) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := iread1_2667(7 downto 0);
      ival1_2735 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2738_inst
    process(iread2_2676) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := iread2_2676(7 downto 0);
      ival2_2739 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2742_inst
    process(iread3_2685) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := iread3_2685(7 downto 0);
      ival3_2743 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2746_inst
    process(iread4_2694) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := iread4_2694(7 downto 0);
      ival4_2747 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2810_inst
    process(kread1_2789) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kread1_2789(7 downto 0);
      kval1_2811 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2814_inst
    process(kread2_2798) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kread2_2798(7 downto 0);
      kval2_2815 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2818_inst
    process(kread3_2807) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kread3_2807(7 downto 0);
      kval3_2819 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2824_inst
    process(MUL_i8_i8_2823_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2823_wire(7 downto 0);
      mul_val1_2825 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2830_inst
    process(MUL_i8_i8_2829_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2829_wire(7 downto 0);
      mul_val2_2831 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2836_inst
    process(MUL_i8_i8_2835_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2835_wire(7 downto 0);
      mul_val3_2837 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2842_inst
    process(MUL_i8_i8_2841_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2841_wire(7 downto 0);
      mul_val4_2843 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2848_inst
    process(MUL_i8_i8_2847_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2847_wire(7 downto 0);
      mul_val5_2849 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2854_inst
    process(MUL_i8_i8_2853_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2853_wire(7 downto 0);
      mul_val6_2855 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3006_inst
    process(acc_val1_2867) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := acc_val1_2867(7 downto 0);
      type_cast_3006_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3008_inst
    process(acc_val2_2879) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := acc_val2_2879(7 downto 0);
      type_cast_3008_wire <= tmp_var; -- 
    end process;
    do_while_stmt_2583_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_3013_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2583_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2583_branch_req_0,
          ack0 => do_while_stmt_2583_branch_ack_0,
          ack1 => do_while_stmt_2583_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i8_i8_2862_inst
    process(acc1_2767_delayed_1_0_2858, mul_val1_2825) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(acc1_2767_delayed_1_0_2858, mul_val1_2825, tmp_var);
      ADD_i8_i8_2862_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2865_inst
    process(mul_val2_2831, mul_val3_2837) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val2_2831, mul_val3_2837, tmp_var);
      ADD_i8_i8_2865_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2866_inst
    process(ADD_i8_i8_2862_wire, ADD_i8_i8_2865_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2862_wire, ADD_i8_i8_2865_wire, tmp_var);
      acc_val1_2867 <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2874_inst
    process(acc2_2776_delayed_1_0_2870, mul_val4_2843) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(acc2_2776_delayed_1_0_2870, mul_val4_2843, tmp_var);
      ADD_i8_i8_2874_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2877_inst
    process(mul_val5_2849, mul_val6_2855) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val5_2849, mul_val6_2855, tmp_var);
      ADD_i8_i8_2877_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2878_inst
    process(ADD_i8_i8_2874_wire, ADD_i8_i8_2877_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2874_wire, ADD_i8_i8_2877_wire, tmp_var);
      acc_val2_2879 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2949_inst
    process(chl_2612) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_2612, konst_2948_wire_constant, tmp_var);
      ADD_u16_u16_2949_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2969_inst
    process(col_2601) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_2601, konst_2968_wire_constant, tmp_var);
      ADD_u16_u16_2969_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2978_inst
    process(row_2596) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_2596, konst_2977_wire_constant, tmp_var);
      ADD_u16_u16_2978_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u2_u2_2958_inst
    process(num_2606) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_2606, konst_2957_wire_constant, tmp_var);
      ADD_u2_u2_2958_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2702_inst
    process(ULT_u16_u1_2698_wire, UGT_u2_u1_2701_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ULT_u16_u1_2698_wire, UGT_u2_u1_2701_wire, tmp_var);
      write_input_2703 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2755_inst
    process(EQ_u16_u1_2751_wire, EQ_u16_u1_2754_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u16_u1_2751_wire, EQ_u16_u1_2754_wire, tmp_var);
      read_k_2756 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2890_inst
    process(EQ_u2_u1_2888_wire, chl_done_2884) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_2888_wire, chl_done_2884, tmp_var);
      num_done_2891 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2900_inst
    process(col_done_2896, num_done_2891) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_2896, num_done_2891, tmp_var);
      row_done_2901 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2915_inst
    process(out_done_flag_2911, col_done_2896) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_2911, col_done_2896, tmp_var);
      AND_u1_u1_2915_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2921_inst
    process(out_done_flag_2911, row_done_2901) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_2911, row_done_2901, tmp_var);
      all_done_flag_2922 <= tmp_var; --
    end process;
    -- shared split operator group (16) : CONCAT_u8_u16_3009_inst 
    ApConcat_group_16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3006_wire & type_cast_3008_wire;
      CONCAT_u8_u16_3009_wire <= data_out(15 downto 0);
      guard_vector(0)  <= num_done_2886_delayed_1_0_3002(0);
      reqL_unguarded(0) <= CONCAT_u8_u16_3009_inst_req_0;
      CONCAT_u8_u16_3009_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u8_u16_3009_inst_req_1;
      CONCAT_u8_u16_3009_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_16_gI: SplitGuardInterface generic map(name => "ApConcat_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- binary operator EQ_u16_u1_2621_inst
    process(col_2601) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2601, konst_2620_wire_constant, tmp_var);
      EQ_u16_u1_2621_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2751_inst
    process(col_2601) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2601, konst_2750_wire_constant, tmp_var);
      EQ_u16_u1_2751_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2754_inst
    process(row_2596) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(row_2596, konst_2753_wire_constant, tmp_var);
      EQ_u16_u1_2754_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2883_inst
    process(chl_2612, num_chl_2582) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(chl_2612, num_chl_2582, tmp_var);
      chl_done_2884 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2895_inst
    process(col_2601, num_col_2577) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2601, num_col_2577, tmp_var);
      col_done_2896 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2624_inst
    process(num_2606) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_2606, konst_2623_wire_constant, tmp_var);
      EQ_u2_u1_2624_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2888_inst
    process(num_2606) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_2606, konst_2887_wire_constant, tmp_var);
      EQ_u2_u1_2888_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2823_inst
    process(kval1_2811, ival1_2735) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_2811, ival1_2735, tmp_var);
      MUL_i8_i8_2823_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2829_inst
    process(kval2_2815, ival2_2739) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_2815, ival2_2739, tmp_var);
      MUL_i8_i8_2829_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2835_inst
    process(kval3_2819, ival3_2743) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_2819, ival3_2743, tmp_var);
      MUL_i8_i8_2835_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2841_inst
    process(kval1_2811, ival2_2739) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_2811, ival2_2739, tmp_var);
      MUL_i8_i8_2841_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2847_inst
    process(kval2_2815, ival3_2743) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_2815, ival3_2743, tmp_var);
      MUL_i8_i8_2847_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2853_inst
    process(kval3_2819, ival4_2747) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_2819, ival4_2747, tmp_var);
      MUL_i8_i8_2853_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2916_inst
    process(AND_u1_u1_2915_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", AND_u1_u1_2915_wire, tmp_var);
      store_kernel_2917 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3013_inst
    process(all_done_flag_2922) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", all_done_flag_2922, tmp_var);
      NOT_u1_u1_3013_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2625_inst
    process(EQ_u16_u1_2621_wire, EQ_u2_u1_2624_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u16_u1_2621_wire, EQ_u2_u1_2624_wire, tmp_var);
      read_ip_2626 <= tmp_var; --
    end process;
    -- shared split operator group (33) : SUB_u16_u16_2571_inst 
    ApIntSub_group_33: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_2569_wire;
      num_row_2572 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2571_inst_req_0;
      SUB_u16_u16_2571_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2571_inst_req_1;
      SUB_u16_u16_2571_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_33_gI: SplitGuardInterface generic map(name => "ApIntSub_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : SUB_u16_u16_2576_inst 
    ApIntSub_group_34: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_2574_wire;
      num_col_2577 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2576_inst_req_0;
      SUB_u16_u16_2576_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2576_inst_req_1;
      SUB_u16_u16_2576_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_34_gI: SplitGuardInterface generic map(name => "ApIntSub_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : SUB_u16_u16_2581_inst 
    ApIntSub_group_35: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_size_pipe_2579_wire;
      num_chl_2582 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2581_inst_req_0;
      SUB_u16_u16_2581_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2581_inst_req_1;
      SUB_u16_u16_2581_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_35_gI: SplitGuardInterface generic map(name => "ApIntSub_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : SUB_u16_u16_2905_inst 
    ApIntSub_group_36: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= num_row_2572;
      SUB_u16_u16_2810_2810_delayed_1_0_2906 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2905_inst_req_0;
      SUB_u16_u16_2905_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2905_inst_req_1;
      SUB_u16_u16_2905_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_36_gI: SplitGuardInterface generic map(name => "ApIntSub_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- binary operator UGE_u16_u1_2910_inst
    process(row_2596, SUB_u16_u16_2810_2810_delayed_1_0_2906) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(row_2596, SUB_u16_u16_2810_2810_delayed_1_0_2906, tmp_var);
      out_done_flag_2911 <= tmp_var; --
    end process;
    -- binary operator UGT_u2_u1_2701_inst
    process(num_2606) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_2606, konst_2700_wire_constant, tmp_var);
      UGT_u2_u1_2701_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_2698_inst
    process(col_2601, num_col_2577) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(col_2601, num_col_2577, tmp_var);
      ULT_u16_u1_2698_wire <= tmp_var; --
    end process;
    xxconvolvexxconv_ip1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip1",
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip1_pipe_read_req,
        read_ack => xxconvolvexxconv_ip1_pipe_read_ack,
        read_data => xxconvolvexxconv_ip1_pipe_read_data,
        write_req => xxconvolvexxconv_ip1_pipe_write_req,
        write_ack => xxconvolvexxconv_ip1_pipe_write_ack,
        write_data => xxconvolvexxconv_ip1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip2",
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip2_pipe_read_req,
        read_ack => xxconvolvexxconv_ip2_pipe_read_ack,
        read_data => xxconvolvexxconv_ip2_pipe_read_data,
        write_req => xxconvolvexxconv_ip2_pipe_write_req,
        write_ack => xxconvolvexxconv_ip2_pipe_write_ack,
        write_data => xxconvolvexxconv_ip2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip3",
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip3_pipe_read_req,
        read_ack => xxconvolvexxconv_ip3_pipe_read_ack,
        read_data => xxconvolvexxconv_ip3_pipe_read_data,
        write_req => xxconvolvexxconv_ip3_pipe_write_req,
        write_ack => xxconvolvexxconv_ip3_pipe_write_ack,
        write_data => xxconvolvexxconv_ip3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip4_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip4",
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip4_pipe_read_req,
        read_ack => xxconvolvexxconv_ip4_pipe_read_ack,
        read_data => xxconvolvexxconv_ip4_pipe_read_data,
        write_req => xxconvolvexxconv_ip4_pipe_write_req,
        write_ack => xxconvolvexxconv_ip4_pipe_write_ack,
        write_data => xxconvolvexxconv_ip4_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k1",
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k1_pipe_read_req,
        read_ack => xxconvolvexxconv_k1_pipe_read_ack,
        read_data => xxconvolvexxconv_k1_pipe_read_data,
        write_req => xxconvolvexxconv_k1_pipe_write_req,
        write_ack => xxconvolvexxconv_k1_pipe_write_ack,
        write_data => xxconvolvexxconv_k1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k2",
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k2_pipe_read_req,
        read_ack => xxconvolvexxconv_k2_pipe_read_ack,
        read_data => xxconvolvexxconv_k2_pipe_read_data,
        write_req => xxconvolvexxconv_k2_pipe_write_req,
        write_ack => xxconvolvexxconv_k2_pipe_write_ack,
        write_data => xxconvolvexxconv_k2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k3",
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k3_pipe_read_req,
        read_ack => xxconvolvexxconv_k3_pipe_read_ack,
        read_data => xxconvolvexxconv_k3_pipe_read_data,
        write_req => xxconvolvexxconv_k3_pipe_write_req,
        write_ack => xxconvolvexxconv_k3_pipe_write_ack,
        write_data => xxconvolvexxconv_k3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    -- shared inport operator group (0) : RPIPE_input_pipe1_2629_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_2629_inst_req_0;
      RPIPE_input_pipe1_2629_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_2629_inst_req_1;
      RPIPE_input_pipe1_2629_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2626(0);
      temp2_1_2630 <= data_out(7 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_input_pipe2_2633_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe2_2633_inst_req_0;
      RPIPE_input_pipe2_2633_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe2_2633_inst_req_1;
      RPIPE_input_pipe2_2633_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2626(0);
      temp2_2_2634 <= data_out(7 downto 0);
      input_pipe2_read_1_gI: SplitGuardInterface generic map(name => "input_pipe2_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe2_read_1: InputPortRevised -- 
        generic map ( name => "input_pipe2_read_1", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe2_pipe_read_req(0),
          oack => input_pipe2_pipe_read_ack(0),
          odata => input_pipe2_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_input_pipe3_2637_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe3_2637_inst_req_0;
      RPIPE_input_pipe3_2637_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe3_2637_inst_req_1;
      RPIPE_input_pipe3_2637_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2626(0);
      temp2_3_2638 <= data_out(7 downto 0);
      input_pipe3_read_2_gI: SplitGuardInterface generic map(name => "input_pipe3_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe3_read_2: InputPortRevised -- 
        generic map ( name => "input_pipe3_read_2", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe3_pipe_read_req(0),
          oack => input_pipe3_pipe_read_ack(0),
          odata => input_pipe3_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_input_pipe4_2641_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe4_2641_inst_req_0;
      RPIPE_input_pipe4_2641_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe4_2641_inst_req_1;
      RPIPE_input_pipe4_2641_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2626(0);
      temp2_4_2642 <= data_out(7 downto 0);
      input_pipe4_read_3_gI: SplitGuardInterface generic map(name => "input_pipe4_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe4_read_3: InputPortRevised -- 
        generic map ( name => "input_pipe4_read_3", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe4_pipe_read_req(0),
          oack => input_pipe4_pipe_read_ack(0),
          odata => input_pipe4_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_kernel_pipe1_2759_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_2759_inst_req_0;
      RPIPE_kernel_pipe1_2759_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_2759_inst_req_1;
      RPIPE_kernel_pipe1_2759_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2756(0);
      tempk1_1_2760 <= data_out(7 downto 0);
      kernel_pipe1_read_4_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_4: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_4", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : RPIPE_kernel_pipe2_2763_inst 
    InportGroup_5: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe2_2763_inst_req_0;
      RPIPE_kernel_pipe2_2763_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe2_2763_inst_req_1;
      RPIPE_kernel_pipe2_2763_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2756(0);
      tempk1_2_2764 <= data_out(7 downto 0);
      kernel_pipe2_read_5_gI: SplitGuardInterface generic map(name => "kernel_pipe2_read_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_read_5: InputPortRevised -- 
        generic map ( name => "kernel_pipe2_read_5", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe2_pipe_read_req(0),
          oack => kernel_pipe2_pipe_read_ack(0),
          odata => kernel_pipe2_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : RPIPE_kernel_pipe3_2767_inst 
    InportGroup_6: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe3_2767_inst_req_0;
      RPIPE_kernel_pipe3_2767_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe3_2767_inst_req_1;
      RPIPE_kernel_pipe3_2767_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2756(0);
      tempk1_3_2768 <= data_out(7 downto 0);
      kernel_pipe3_read_6_gI: SplitGuardInterface generic map(name => "kernel_pipe3_read_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_read_6: InputPortRevised -- 
        generic map ( name => "kernel_pipe3_read_6", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe3_pipe_read_req(0),
          oack => kernel_pipe3_pipe_read_ack(0),
          odata => kernel_pipe3_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : RPIPE_num_out_pipe_2569_inst RPIPE_num_out_pipe_2574_inst 
    InportGroup_7: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_num_out_pipe_2569_inst_req_0;
      reqL_unguarded(0) <= RPIPE_num_out_pipe_2574_inst_req_0;
      RPIPE_num_out_pipe_2569_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_num_out_pipe_2574_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_num_out_pipe_2569_inst_req_1;
      reqR_unguarded(0) <= RPIPE_num_out_pipe_2574_inst_req_1;
      RPIPE_num_out_pipe_2569_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_num_out_pipe_2574_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      RPIPE_num_out_pipe_2569_wire <= data_out(31 downto 16);
      RPIPE_num_out_pipe_2574_wire <= data_out(15 downto 0);
      num_out_pipe_read_7_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_7_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_7: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_7", data_width => 16,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : RPIPE_size_pipe_2579_inst 
    InportGroup_8: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_2579_inst_req_0;
      RPIPE_size_pipe_2579_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_2579_inst_req_1;
      RPIPE_size_pipe_2579_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_size_pipe_2579_wire <= data_out(15 downto 0);
      size_pipe_read_8_gI: SplitGuardInterface generic map(name => "size_pipe_read_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_8: InputPortRevised -- 
        generic map ( name => "size_pipe_read_8", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared inport operator group (9) : RPIPE_xxconvolvexxconv_ip1_2645_inst 
    InportGroup_9: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_2645_inst_req_0;
      RPIPE_xxconvolvexxconv_ip1_2645_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_2645_inst_req_1;
      RPIPE_xxconvolvexxconv_ip1_2645_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2626(0);
      temp1_1_2646 <= data_out(7 downto 0);
      xxconvolvexxconv_ip1_read_9_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_read_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_read_9: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1_read_9", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip1_pipe_read_req(0),
          oack => xxconvolvexxconv_ip1_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 9
    -- shared inport operator group (10) : RPIPE_xxconvolvexxconv_ip2_2649_inst 
    InportGroup_10: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_2649_inst_req_0;
      RPIPE_xxconvolvexxconv_ip2_2649_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_2649_inst_req_1;
      RPIPE_xxconvolvexxconv_ip2_2649_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2626(0);
      temp1_2_2650 <= data_out(7 downto 0);
      xxconvolvexxconv_ip2_read_10_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_read_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_read_10: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2_read_10", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip2_pipe_read_req(0),
          oack => xxconvolvexxconv_ip2_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 10
    -- shared inport operator group (11) : RPIPE_xxconvolvexxconv_ip3_2653_inst 
    InportGroup_11: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_2653_inst_req_0;
      RPIPE_xxconvolvexxconv_ip3_2653_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_2653_inst_req_1;
      RPIPE_xxconvolvexxconv_ip3_2653_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2626(0);
      temp1_3_2654 <= data_out(7 downto 0);
      xxconvolvexxconv_ip3_read_11_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_read_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_read_11: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3_read_11", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip3_pipe_read_req(0),
          oack => xxconvolvexxconv_ip3_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 11
    -- shared inport operator group (12) : RPIPE_xxconvolvexxconv_ip4_2657_inst 
    InportGroup_12: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip4_2657_inst_req_0;
      RPIPE_xxconvolvexxconv_ip4_2657_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip4_2657_inst_req_1;
      RPIPE_xxconvolvexxconv_ip4_2657_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2626(0);
      temp1_4_2658 <= data_out(7 downto 0);
      xxconvolvexxconv_ip4_read_12_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip4_read_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip4_read_12: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip4_read_12", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip4_pipe_read_req(0),
          oack => xxconvolvexxconv_ip4_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip4_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 12
    -- shared inport operator group (13) : RPIPE_xxconvolvexxconv_k1_2771_inst 
    InportGroup_13: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_2771_inst_req_0;
      RPIPE_xxconvolvexxconv_k1_2771_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_2771_inst_req_1;
      RPIPE_xxconvolvexxconv_k1_2771_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2756(0);
      tempk2_1_2772 <= data_out(7 downto 0);
      xxconvolvexxconv_k1_read_13_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_read_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_read_13: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1_read_13", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k1_pipe_read_req(0),
          oack => xxconvolvexxconv_k1_pipe_read_ack(0),
          odata => xxconvolvexxconv_k1_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 13
    -- shared inport operator group (14) : RPIPE_xxconvolvexxconv_k2_2775_inst 
    InportGroup_14: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_2775_inst_req_0;
      RPIPE_xxconvolvexxconv_k2_2775_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_2775_inst_req_1;
      RPIPE_xxconvolvexxconv_k2_2775_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2756(0);
      tempk2_2_2776 <= data_out(7 downto 0);
      xxconvolvexxconv_k2_read_14_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_read_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_read_14: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2_read_14", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k2_pipe_read_req(0),
          oack => xxconvolvexxconv_k2_pipe_read_ack(0),
          odata => xxconvolvexxconv_k2_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 14
    -- shared inport operator group (15) : RPIPE_xxconvolvexxconv_k3_2779_inst 
    InportGroup_15: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_2779_inst_req_0;
      RPIPE_xxconvolvexxconv_k3_2779_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_2779_inst_req_1;
      RPIPE_xxconvolvexxconv_k3_2779_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2756(0);
      tempk2_3_2780 <= data_out(7 downto 0);
      xxconvolvexxconv_k3_read_15_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_read_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_read_15: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3_read_15", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k3_pipe_read_req(0),
          oack => xxconvolvexxconv_k3_pipe_read_ack(0),
          odata => xxconvolvexxconv_k3_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 15
    -- shared outport operator group (0) : WPIPE_input_done_pipe_3014_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_3014_inst_req_0;
      WPIPE_input_done_pipe_3014_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_3014_inst_req_1;
      WPIPE_input_done_pipe_3014_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_3015_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_output_pipe_3004_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_output_pipe_3004_inst_req_0;
      WPIPE_output_pipe_3004_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_output_pipe_3004_inst_req_1;
      WPIPE_output_pipe_3004_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= num_done_2886_delayed_1_0_3002(0);
      data_in <= CONCAT_u8_u16_3009_wire;
      output_pipe_write_1_gI: SplitGuardInterface generic map(name => "output_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "output_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => output_pipe_pipe_write_req(0),
          oack => output_pipe_pipe_write_ack(0),
          odata => output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_xxconvolvexxconv_ip1_2708_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_2708_inst_req_0;
      WPIPE_xxconvolvexxconv_ip1_2708_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_2708_inst_req_1;
      WPIPE_xxconvolvexxconv_ip1_2708_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2635_delayed_1_0_2706(0);
      data_in <= iread1_2667;
      xxconvolvexxconv_ip1_write_2_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_write_2: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip1_pipe_write_req(0),
          oack => xxconvolvexxconv_ip1_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_xxconvolvexxconv_ip2_2715_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_2715_inst_req_0;
      WPIPE_xxconvolvexxconv_ip2_2715_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_2715_inst_req_1;
      WPIPE_xxconvolvexxconv_ip2_2715_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2639_delayed_1_0_2713(0);
      data_in <= iread2_2676;
      xxconvolvexxconv_ip2_write_3_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_write_3: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip2_pipe_write_req(0),
          oack => xxconvolvexxconv_ip2_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_xxconvolvexxconv_ip3_2722_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_2722_inst_req_0;
      WPIPE_xxconvolvexxconv_ip3_2722_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_2722_inst_req_1;
      WPIPE_xxconvolvexxconv_ip3_2722_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2643_delayed_1_0_2720(0);
      data_in <= iread3_2685;
      xxconvolvexxconv_ip3_write_4_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_write_4: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip3_pipe_write_req(0),
          oack => xxconvolvexxconv_ip3_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_xxconvolvexxconv_ip4_2729_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip4_2729_inst_req_0;
      WPIPE_xxconvolvexxconv_ip4_2729_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip4_2729_inst_req_1;
      WPIPE_xxconvolvexxconv_ip4_2729_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2647_delayed_1_0_2727(0);
      data_in <= iread4_2694;
      xxconvolvexxconv_ip4_write_5_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip4_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip4_write_5: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip4", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip4_pipe_write_req(0),
          oack => xxconvolvexxconv_ip4_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip4_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared outport operator group (6) : WPIPE_xxconvolvexxconv_k1_2927_inst 
    OutportGroup_6: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_2927_inst_req_0;
      WPIPE_xxconvolvexxconv_k1_2927_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_2927_inst_req_1;
      WPIPE_xxconvolvexxconv_k1_2927_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2824_delayed_1_0_2925(0);
      data_in <= kread1_2789;
      xxconvolvexxconv_k1_write_6_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_write_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_write_6: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k1_pipe_write_req(0),
          oack => xxconvolvexxconv_k1_pipe_write_ack(0),
          odata => xxconvolvexxconv_k1_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- shared outport operator group (7) : WPIPE_xxconvolvexxconv_k2_2934_inst 
    OutportGroup_7: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_2934_inst_req_0;
      WPIPE_xxconvolvexxconv_k2_2934_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_2934_inst_req_1;
      WPIPE_xxconvolvexxconv_k2_2934_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2828_delayed_1_0_2932(0);
      data_in <= kread2_2798;
      xxconvolvexxconv_k2_write_7_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_write_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_write_7: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k2_pipe_write_req(0),
          oack => xxconvolvexxconv_k2_pipe_write_ack(0),
          odata => xxconvolvexxconv_k2_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- shared outport operator group (8) : WPIPE_xxconvolvexxconv_k3_2941_inst 
    OutportGroup_8: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_2941_inst_req_0;
      WPIPE_xxconvolvexxconv_k3_2941_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_2941_inst_req_1;
      WPIPE_xxconvolvexxconv_k3_2941_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2832_delayed_1_0_2939(0);
      data_in <= kread3_2807;
      xxconvolvexxconv_k3_write_8_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_write_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_write_8: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k3_pipe_write_req(0),
          oack => xxconvolvexxconv_k3_pipe_write_ack(0),
          odata => xxconvolvexxconv_k3_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 8
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    num_chl : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_data : out  std_logic_vector(7 downto 0);
    kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_data : out  std_logic_vector(7 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(7 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal num_chl_buffer :  std_logic_vector(15 downto 0);
  signal num_chl_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_1635_start: Boolean;
  signal loadKernelChannel_CP_1635_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nmycount_603_584_buf_ack_1 : boolean;
  signal RPIPE_input_done_pipe_576_inst_ack_1 : boolean;
  signal addr_of_543_final_reg_req_0 : boolean;
  signal RPIPE_input_done_pipe_576_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_576_inst_ack_0 : boolean;
  signal addr_of_543_final_reg_ack_0 : boolean;
  signal nmycount_603_584_buf_req_0 : boolean;
  signal my_fetch_548_588_buf_req_1 : boolean;
  signal nmycount_603_584_buf_ack_0 : boolean;
  signal array_obj_ref_542_index_offset_ack_1 : boolean;
  signal ptr_deref_547_load_0_ack_0 : boolean;
  signal ptr_deref_547_load_0_req_0 : boolean;
  signal array_obj_ref_542_index_offset_req_1 : boolean;
  signal ptr_deref_547_load_0_ack_1 : boolean;
  signal RPIPE_input_done_pipe_576_inst_req_1 : boolean;
  signal ptr_deref_547_load_0_req_1 : boolean;
  signal start_add_583_buf_ack_1 : boolean;
  signal array_obj_ref_542_index_offset_ack_0 : boolean;
  signal phi_stmt_585_req_1 : boolean;
  signal array_obj_ref_542_index_offset_req_0 : boolean;
  signal nfetch_val_675_587_buf_ack_0 : boolean;
  signal start_add_583_buf_req_1 : boolean;
  signal nmycount_603_584_buf_req_1 : boolean;
  signal nfetch_val_675_587_buf_req_0 : boolean;
  signal phi_stmt_585_ack_0 : boolean;
  signal nfetch_val_675_587_buf_req_1 : boolean;
  signal nfetch_val_675_587_buf_ack_1 : boolean;
  signal my_fetch_548_588_buf_req_0 : boolean;
  signal phi_stmt_581_req_1 : boolean;
  signal addr_of_543_final_reg_req_1 : boolean;
  signal my_fetch_548_588_buf_ack_1 : boolean;
  signal addr_of_543_final_reg_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_629_inst_ack_1 : boolean;
  signal start_add_583_buf_req_0 : boolean;
  signal my_fetch_548_588_buf_ack_0 : boolean;
  signal start_add_583_buf_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_629_inst_req_0 : boolean;
  signal phi_stmt_585_req_0 : boolean;
  signal do_while_stmt_579_branch_req_0 : boolean;
  signal phi_stmt_581_req_0 : boolean;
  signal WPIPE_kernel_pipe1_629_inst_req_1 : boolean;
  signal array_obj_ref_653_index_offset_req_0 : boolean;
  signal phi_stmt_581_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_633_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_633_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe3_637_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe3_637_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe3_637_inst_ack_1 : boolean;
  signal array_obj_ref_653_index_offset_ack_0 : boolean;
  signal array_obj_ref_653_index_offset_req_1 : boolean;
  signal array_obj_ref_653_index_offset_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_629_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_633_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe2_633_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe3_637_inst_req_0 : boolean;
  signal addr_of_654_final_reg_req_0 : boolean;
  signal addr_of_654_final_reg_ack_0 : boolean;
  signal addr_of_654_final_reg_req_1 : boolean;
  signal addr_of_654_final_reg_ack_1 : boolean;
  signal W_fn_608_delayed_7_0_656_inst_req_0 : boolean;
  signal W_fn_608_delayed_7_0_656_inst_ack_0 : boolean;
  signal W_fn_608_delayed_7_0_656_inst_req_1 : boolean;
  signal W_fn_608_delayed_7_0_656_inst_ack_1 : boolean;
  signal ptr_deref_662_load_0_req_0 : boolean;
  signal ptr_deref_662_load_0_ack_0 : boolean;
  signal ptr_deref_662_load_0_req_1 : boolean;
  signal ptr_deref_662_load_0_ack_1 : boolean;
  signal W_fn_614_delayed_13_0_664_inst_req_0 : boolean;
  signal W_fn_614_delayed_13_0_664_inst_ack_0 : boolean;
  signal W_fn_614_delayed_13_0_664_inst_req_1 : boolean;
  signal W_fn_614_delayed_13_0_664_inst_ack_1 : boolean;
  signal W_fetch_val_616_delayed_13_0_667_inst_req_0 : boolean;
  signal W_fetch_val_616_delayed_13_0_667_inst_ack_0 : boolean;
  signal W_fetch_val_616_delayed_13_0_667_inst_req_1 : boolean;
  signal W_fetch_val_616_delayed_13_0_667_inst_ack_1 : boolean;
  signal do_while_stmt_579_branch_ack_0 : boolean;
  signal do_while_stmt_579_branch_ack_1 : boolean;
  signal WPIPE_size_pipe_683_inst_req_0 : boolean;
  signal WPIPE_size_pipe_683_inst_ack_0 : boolean;
  signal WPIPE_size_pipe_683_inst_req_1 : boolean;
  signal WPIPE_size_pipe_683_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(79 downto 64) <= num_chl;
  num_chl_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_1635_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1635_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1635_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1635_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_1635: Block -- control-path 
    signal loadKernelChannel_CP_1635_elements: BooleanArray(98 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_1635_elements(0) <= loadKernelChannel_CP_1635_start;
    loadKernelChannel_CP_1635_symbol <= loadKernelChannel_CP_1635_elements(98);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_complete/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_sample_start_
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Sample/rr
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_complete/req
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_update_start
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_update_start_
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_computed_1
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_resized_1
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_update_start_
      -- 
    req_1685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(0), ack => addr_of_543_final_reg_req_1); -- 
    req_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(0), ack => array_obj_ref_542_index_offset_req_0); -- 
    req_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(0), ack => array_obj_ref_542_index_offset_req_1); -- 
    cr_1730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(0), ack => ptr_deref_547_load_0_req_1); -- 
    rr_1744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(0), ack => RPIPE_input_done_pipe_576_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Sample/ack
      -- CP-element group 1: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_sample_complete
      -- 
    ack_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_542_index_offset_ack_0, ack => loadKernelChannel_CP_1635_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_request/req
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_request/$entry
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_sample_start_
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_offset_calculated
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_root_address_calculated
      -- 
    ack_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_542_index_offset_ack_1, ack => loadKernelChannel_CP_1635_elements(2)); -- 
    req_1680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(2), ack => addr_of_543_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_request/$exit
      -- CP-element group 3: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_request/ack
      -- CP-element group 3: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_sample_completed_
      -- 
    ack_1681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_543_final_reg_ack_0, ack => loadKernelChannel_CP_1635_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_address_resized
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_complete/$exit
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/word_0/rr
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_complete/ack
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_sample_start_
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_update_completed_
      -- 
    ack_1686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_543_final_reg_ack_1, ack => loadKernelChannel_CP_1635_elements(4)); -- 
    rr_1719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(4), ack => ptr_deref_547_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_sample_completed_
      -- CP-element group 5: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/$exit
      -- 
    ra_1720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_547_load_0_ack_0, ack => loadKernelChannel_CP_1635_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/ptr_deref_547_Merge/merge_ack
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/ptr_deref_547_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/ptr_deref_547_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/ptr_deref_547_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/$exit
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_update_completed_
      -- 
    ca_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_547_load_0_ack_1, ack => loadKernelChannel_CP_1635_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_update_start_
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_sample_completed_
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Sample/ra
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Update/$entry
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Update/cr
      -- 
    ra_1745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_576_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(7)); -- 
    cr_1749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(7), ack => RPIPE_input_done_pipe_576_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Update/ca
      -- CP-element group 8: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_update_completed_
      -- CP-element group 8: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Update/$exit
      -- 
    ca_1750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_576_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_578/do_while_stmt_579__entry__
      -- CP-element group 9: 	 branch_block_stmt_578/$entry
      -- CP-element group 9: 	 branch_block_stmt_578/branch_block_stmt_578__entry__
      -- CP-element group 9: 	 assign_stmt_532_to_assign_stmt_577/$exit
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(1) & loadKernelChannel_CP_1635_elements(6) & loadKernelChannel_CP_1635_elements(8);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	96 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	97 
    -- CP-element group 10:  members (7) 
      -- CP-element group 10: 	 branch_block_stmt_578/branch_block_stmt_578__exit__
      -- CP-element group 10: 	 branch_block_stmt_578/do_while_stmt_579__exit__
      -- CP-element group 10: 	 branch_block_stmt_578/$exit
      -- CP-element group 10: 	 assign_stmt_685/$entry
      -- CP-element group 10: 	 assign_stmt_685/WPIPE_size_pipe_683_sample_start_
      -- CP-element group 10: 	 assign_stmt_685/WPIPE_size_pipe_683_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_685/WPIPE_size_pipe_683_Sample/req
      -- 
    req_2086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(10), ack => WPIPE_size_pipe_683_inst_req_0); -- 
    loadKernelChannel_CP_1635_elements(10) <= loadKernelChannel_CP_1635_elements(96);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579__entry__
      -- CP-element group 11: 	 branch_block_stmt_578/do_while_stmt_579/$entry
      -- 
    loadKernelChannel_CP_1635_elements(11) <= loadKernelChannel_CP_1635_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	96 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579__exit__
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_578/do_while_stmt_579/loop_back
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	94 
    -- CP-element group 14: 	95 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_578/do_while_stmt_579/condition_done
      -- CP-element group 14: 	 branch_block_stmt_578/do_while_stmt_579/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_578/do_while_stmt_579/loop_taken/$entry
      -- 
    loadKernelChannel_CP_1635_elements(14) <= loadKernelChannel_CP_1635_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	93 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_578/do_while_stmt_579/loop_body_done
      -- 
    loadKernelChannel_CP_1635_elements(15) <= loadKernelChannel_CP_1635_elements(93);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	28 
    -- CP-element group 16: 	47 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_1635_elements(16) <= loadKernelChannel_CP_1635_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	49 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_1635_elements(17) <= loadKernelChannel_CP_1635_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	25 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	70 
    -- CP-element group 18: 	71 
    -- CP-element group 18: 	92 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	27 
    -- CP-element group 19: 	92 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/condition_evaluated
      -- 
    condition_evaluated_1772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(19), ack => do_while_stmt_579_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(23) & loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(92);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	41 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	43 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_sample_start__ps
      -- CP-element group 20: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/aggregated_phi_sample_req
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(24) & loadKernelChannel_CP_1635_elements(41) & loadKernelChannel_CP_1635_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: 	44 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	81 
    -- CP-element group 21: 	85 
    -- CP-element group 21: 	89 
    -- CP-element group 21: 	93 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	41 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(26) & loadKernelChannel_CP_1635_elements(44);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	42 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	45 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/aggregated_phi_update_req
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(25) & loadKernelChannel_CP_1635_elements(42);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(46);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	64 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	78 
    -- CP-element group 25: 	86 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(61) & loadKernelChannel_CP_1635_elements(64) & loadKernelChannel_CP_1635_elements(67) & loadKernelChannel_CP_1635_elements(72) & loadKernelChannel_CP_1635_elements(78) & loadKernelChannel_CP_1635_elements(86);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	19 
    -- CP-element group 27: 	23 
    -- CP-element group 27: 	60 
    -- CP-element group 27: 	63 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	72 
    -- CP-element group 27: 	76 
    -- CP-element group 27: 	84 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (15) 
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_scale_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_scale_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_scale_1/scale_rename_req
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_scale_1/scale_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Sample/req
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_resized_1
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_scaled_1
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_computed_1
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_resize_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_resize_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_resize_1/index_resize_req
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_resize_1/index_resize_ack
      -- 
    req_1952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(27), ack => array_obj_ref_653_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	16 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_loopback_trigger
      -- 
    loadKernelChannel_CP_1635_elements(28) <= loadKernelChannel_CP_1635_elements(16);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_loopback_sample_req
      -- CP-element group 29: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_loopback_sample_req_ps
      -- 
    phi_stmt_581_loopback_sample_req_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_581_loopback_sample_req_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(29), ack => phi_stmt_581_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_entry_trigger
      -- 
    loadKernelChannel_CP_1635_elements(30) <= loadKernelChannel_CP_1635_elements(17);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_entry_sample_req
      -- CP-element group 31: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_entry_sample_req_ps
      -- 
    phi_stmt_581_entry_sample_req_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_581_entry_sample_req_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(31), ack => phi_stmt_581_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_phi_mux_ack_ps
      -- CP-element group 32: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_phi_mux_ack
      -- 
    phi_stmt_581_phi_mux_ack_1793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_581_ack_0, ack => loadKernelChannel_CP_1635_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Sample/req
      -- 
    req_1806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(33), ack => start_add_583_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_update_start_
      -- CP-element group 34: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Update/req
      -- CP-element group 34: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Update/$entry
      -- 
    req_1811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(34), ack => start_add_583_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Sample/ack
      -- 
    ack_1807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_583_buf_ack_0, ack => loadKernelChannel_CP_1635_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Update/ack
      -- CP-element group 36: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_update_completed__ps
      -- 
    ack_1812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_583_buf_ack_1, ack => loadKernelChannel_CP_1635_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_sample_start__ps
      -- 
    req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(37), ack => nmycount_603_584_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_update_start_
      -- CP-element group 38: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Update/req
      -- CP-element group 38: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_update_start__ps
      -- 
    req_1829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(38), ack => nmycount_603_584_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_sample_completed__ps
      -- 
    ack_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_603_584_buf_ack_0, ack => loadKernelChannel_CP_1635_elements(39)); -- 
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_update_completed__ps
      -- 
    ack_1830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_603_584_buf_ack_1, ack => loadKernelChannel_CP_1635_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	21 
    -- CP-element group 41: 	83 
    -- CP-element group 41: 	87 
    -- CP-element group 41: 	91 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	20 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_sample_start_
      -- 
    loadKernelChannel_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(21) & loadKernelChannel_CP_1635_elements(83) & loadKernelChannel_CP_1635_elements(87) & loadKernelChannel_CP_1635_elements(91);
      gj_loadKernelChannel_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	18 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	46 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	64 
    -- CP-element group 42: 	67 
    -- CP-element group 42: 	90 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	22 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_update_start_
      -- 
    loadKernelChannel_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(46) & loadKernelChannel_CP_1635_elements(61) & loadKernelChannel_CP_1635_elements(64) & loadKernelChannel_CP_1635_elements(67) & loadKernelChannel_CP_1635_elements(90);
      gj_loadKernelChannel_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	20 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_sample_start__ps
      -- 
    loadKernelChannel_CP_1635_elements(43) <= loadKernelChannel_CP_1635_elements(20);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	22 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_update_start__ps
      -- 
    loadKernelChannel_CP_1635_elements(45) <= loadKernelChannel_CP_1635_elements(22);
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	63 
    -- CP-element group 46: 	66 
    -- CP-element group 46: 	88 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	42 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_update_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_update_completed_
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_loopback_trigger
      -- 
    loadKernelChannel_CP_1635_elements(47) <= loadKernelChannel_CP_1635_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_loopback_sample_req
      -- CP-element group 48: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_loopback_sample_req_ps
      -- 
    phi_stmt_585_loopback_sample_req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_585_loopback_sample_req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(48), ack => phi_stmt_585_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_entry_trigger
      -- 
    loadKernelChannel_CP_1635_elements(49) <= loadKernelChannel_CP_1635_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_entry_sample_req_ps
      -- CP-element group 50: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_entry_sample_req
      -- 
    phi_stmt_585_entry_sample_req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_585_entry_sample_req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(50), ack => phi_stmt_585_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_phi_mux_ack_ps
      -- CP-element group 51: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_phi_mux_ack
      -- 
    phi_stmt_585_phi_mux_ack_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_585_ack_0, ack => loadKernelChannel_CP_1635_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_Sample/$entry
      -- 
    req_1860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(52), ack => nfetch_val_675_587_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_Update/req
      -- CP-element group 53: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_update_start_
      -- 
    req_1865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(53), ack => nfetch_val_675_587_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_Sample/$exit
      -- 
    ack_1861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_675_587_buf_ack_0, ack => loadKernelChannel_CP_1635_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_587_Update/ack
      -- 
    ack_1866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_675_587_buf_ack_1, ack => loadKernelChannel_CP_1635_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_sample_start__ps
      -- 
    req_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(56), ack => my_fetch_548_588_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_Update/req
      -- CP-element group 57: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_update_start_
      -- CP-element group 57: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_update_start__ps
      -- CP-element group 57: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_Update/$entry
      -- 
    req_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(57), ack => my_fetch_548_588_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_sample_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_Sample/$exit
      -- 
    ack_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_548_588_buf_ack_0, ack => loadKernelChannel_CP_1635_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_update_completed__ps
      -- CP-element group 59: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_588_Update/$exit
      -- 
    ack_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_548_588_buf_ack_1, ack => loadKernelChannel_CP_1635_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	27 
    -- CP-element group 60: 	46 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Sample/req
      -- 
    req_1893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(60), ack => WPIPE_kernel_pipe1_629_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(46) & loadKernelChannel_CP_1635_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	25 
    -- CP-element group 61: 	42 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Update/req
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_update_start_
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Sample/$exit
      -- 
    ack_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_629_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(61)); -- 
    req_1898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(61), ack => WPIPE_kernel_pipe1_629_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	93 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_update_completed_
      -- 
    ack_1899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_629_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	27 
    -- CP-element group 63: 	46 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_sample_start_
      -- 
    req_1907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(63), ack => WPIPE_kernel_pipe2_633_inst_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(46) & loadKernelChannel_CP_1635_elements(65);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	25 
    -- CP-element group 64: 	42 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_update_start_
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Update/req
      -- 
    ack_1908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_633_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(64)); -- 
    req_1912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(64), ack => WPIPE_kernel_pipe2_633_inst_req_1); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	93 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Update/ack
      -- 
    ack_1913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_633_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	27 
    -- CP-element group 66: 	46 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Sample/req
      -- 
    req_1921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(66), ack => WPIPE_kernel_pipe3_637_inst_req_0); -- 
    loadKernelChannel_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(46) & loadKernelChannel_CP_1635_elements(68);
      gj_loadKernelChannel_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	42 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Update/req
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_update_start_
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Sample/$exit
      -- 
    ack_1922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_637_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(67)); -- 
    req_1926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(67), ack => WPIPE_kernel_pipe3_637_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	93 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_update_completed_
      -- 
    ack_1927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_637_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	73 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_request/$entry
      -- CP-element group 69: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_request/req
      -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(69), ack => addr_of_654_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(73) & loadKernelChannel_CP_1635_elements(74);
      gj_loadKernelChannel_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	18 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	75 
    -- CP-element group 70: 	82 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	75 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_update_start_
      -- CP-element group 70: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_complete/$entry
      -- CP-element group 70: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_complete/req
      -- 
    req_1972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(70), ack => addr_of_654_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(75) & loadKernelChannel_CP_1635_elements(82);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	18 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	74 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_update_start
      -- CP-element group 71: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Update/req
      -- 
    req_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(71), ack => array_obj_ref_653_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(73) & loadKernelChannel_CP_1635_elements(74);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	27 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	93 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	25 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_sample_complete
      -- CP-element group 72: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Sample/ack
      -- 
    ack_1953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_653_index_offset_ack_0, ack => loadKernelChannel_CP_1635_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	69 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (8) 
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_offset_calculated
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_base_plus_offset/sum_rename_ack
      -- 
    ack_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_653_index_offset_ack_1, ack => loadKernelChannel_CP_1635_elements(73)); -- 
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	71 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_request/$exit
      -- CP-element group 74: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_request/ack
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_654_final_reg_ack_0, ack => loadKernelChannel_CP_1635_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	70 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	80 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	70 
    -- CP-element group 75:  members (19) 
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_word_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_complete/ack
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_root_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_address_resized
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_addr_resize/$entry
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_addr_resize/$exit
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_addr_resize/base_resize_req
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_addr_resize/base_resize_ack
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_plus_offset/$entry
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_plus_offset/$exit
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_plus_offset/sum_rename_req
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_plus_offset/sum_rename_ack
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_word_addrgen/$entry
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_word_addrgen/$exit
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_word_addrgen/root_register_req
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_word_addrgen/root_register_ack
      -- 
    ack_1973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_654_final_reg_ack_1, ack => loadKernelChannel_CP_1635_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	27 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Sample/req
      -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(76), ack => W_fn_608_delayed_7_0_656_inst_req_0); -- 
    loadKernelChannel_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(78);
      gj_loadKernelChannel_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	82 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_update_start_
      -- CP-element group 77: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Update/req
      -- 
    req_1986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(77), ack => W_fn_608_delayed_7_0_656_inst_req_1); -- 
    loadKernelChannel_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(79) & loadKernelChannel_CP_1635_elements(82);
      gj_loadKernelChannel_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	25 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Sample/ack
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_608_delayed_7_0_656_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Update/ack
      -- 
    ack_1987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_608_delayed_7_0_656_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: 	79 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/$entry
      -- CP-element group 80: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/word_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/word_0/rr
      -- 
    rr_2020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(80), ack => ptr_deref_662_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(75) & loadKernelChannel_CP_1635_elements(79) & loadKernelChannel_CP_1635_elements(82);
      gj_loadKernelChannel_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	21 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_update_start_
      -- CP-element group 81: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/word_0/cr
      -- 
    cr_2031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(81), ack => ptr_deref_662_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(21) & loadKernelChannel_CP_1635_elements(83);
      gj_loadKernelChannel_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/$exit
      -- CP-element group 82: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/word_0/ra
      -- 
    ra_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_662_load_0_ack_0, ack => loadKernelChannel_CP_1635_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	93 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	41 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/$exit
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/word_0/$exit
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/word_0/ca
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/ptr_deref_662_Merge/$entry
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/ptr_deref_662_Merge/$exit
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/ptr_deref_662_Merge/merge_req
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/ptr_deref_662_Merge/merge_ack
      -- 
    ca_2032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_662_load_0_ack_1, ack => loadKernelChannel_CP_1635_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	27 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Sample/req
      -- 
    req_2045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(84), ack => W_fn_614_delayed_13_0_664_inst_req_0); -- 
    loadKernelChannel_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(86);
      gj_loadKernelChannel_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	21 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_update_start_
      -- CP-element group 85: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Update/req
      -- 
    req_2050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(85), ack => W_fn_614_delayed_13_0_664_inst_req_1); -- 
    loadKernelChannel_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(21) & loadKernelChannel_CP_1635_elements(87);
      gj_loadKernelChannel_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	25 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Sample/ack
      -- 
    ack_2046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_614_delayed_13_0_664_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	93 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	41 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Update/ack
      -- 
    ack_2051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_614_delayed_13_0_664_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	46 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Sample/req
      -- 
    req_2059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(88), ack => W_fetch_val_616_delayed_13_0_667_inst_req_0); -- 
    loadKernelChannel_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(46) & loadKernelChannel_CP_1635_elements(90);
      gj_loadKernelChannel_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	21 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_update_start_
      -- CP-element group 89: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Update/req
      -- 
    req_2064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(89), ack => W_fetch_val_616_delayed_13_0_667_inst_req_1); -- 
    loadKernelChannel_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(21) & loadKernelChannel_CP_1635_elements(91);
      gj_loadKernelChannel_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	42 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Sample/ack
      -- 
    ack_2060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_616_delayed_13_0_667_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	41 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Update/ack
      -- 
    ack_2065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_616_delayed_13_0_667_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(91)); -- 
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	18 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	19 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_1635_elements(18), ack => loadKernelChannel_CP_1635_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	21 
    -- CP-element group 93: 	62 
    -- CP-element group 93: 	65 
    -- CP-element group 93: 	68 
    -- CP-element group 93: 	72 
    -- CP-element group 93: 	83 
    -- CP-element group 93: 	87 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	15 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(21) & loadKernelChannel_CP_1635_elements(62) & loadKernelChannel_CP_1635_elements(65) & loadKernelChannel_CP_1635_elements(68) & loadKernelChannel_CP_1635_elements(72) & loadKernelChannel_CP_1635_elements(83) & loadKernelChannel_CP_1635_elements(87) & loadKernelChannel_CP_1635_elements(91);
      gj_loadKernelChannel_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	14 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_578/do_while_stmt_579/loop_exit/$exit
      -- CP-element group 94: 	 branch_block_stmt_578/do_while_stmt_579/loop_exit/ack
      -- 
    ack_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_579_branch_ack_0, ack => loadKernelChannel_CP_1635_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	14 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_578/do_while_stmt_579/loop_taken/$exit
      -- CP-element group 95: 	 branch_block_stmt_578/do_while_stmt_579/loop_taken/ack
      -- 
    ack_2074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_579_branch_ack_1, ack => loadKernelChannel_CP_1635_elements(95)); -- 
    -- CP-element group 96:  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	12 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	10 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_578/do_while_stmt_579/$exit
      -- 
    loadKernelChannel_CP_1635_elements(96) <= loadKernelChannel_CP_1635_elements(12);
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	10 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_sample_completed_
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_update_start_
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_Sample/$exit
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_Sample/ack
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_Update/$entry
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_Update/req
      -- 
    ack_2087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_683_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(97)); -- 
    req_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(97), ack => WPIPE_size_pipe_683_inst_req_1); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (5) 
      -- CP-element group 98: 	 $exit
      -- CP-element group 98: 	 assign_stmt_685/$exit
      -- CP-element group 98: 	 assign_stmt_685/WPIPE_size_pipe_683_update_completed_
      -- CP-element group 98: 	 assign_stmt_685/WPIPE_size_pipe_683_Update/$exit
      -- CP-element group 98: 	 assign_stmt_685/WPIPE_size_pipe_683_Update/ack
      -- 
    ack_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_683_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(98)); -- 
    loadKernelChannel_do_while_stmt_579_terminator_2075: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_579_terminator_2075", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_1635_elements(15),loop_continue => loadKernelChannel_CP_1635_elements(95),loop_terminate => loadKernelChannel_CP_1635_elements(94),loop_back => loadKernelChannel_CP_1635_elements(13),loop_exit => loadKernelChannel_CP_1635_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_581_phi_seq_1831_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1635_elements(30);
      loadKernelChannel_CP_1635_elements(33)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1635_elements(35);
      loadKernelChannel_CP_1635_elements(34)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1635_elements(36);
      loadKernelChannel_CP_1635_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1635_elements(28);
      loadKernelChannel_CP_1635_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1635_elements(39);
      loadKernelChannel_CP_1635_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1635_elements(40);
      loadKernelChannel_CP_1635_elements(29) <= phi_mux_reqs(1);
      phi_stmt_581_phi_seq_1831 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_581_phi_seq_1831") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1635_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_1635_elements(26), 
          phi_update_req => loadKernelChannel_CP_1635_elements(22), 
          phi_update_ack => loadKernelChannel_CP_1635_elements(27), 
          phi_mux_ack => loadKernelChannel_CP_1635_elements(32), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_585_phi_seq_1885_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1635_elements(47);
      loadKernelChannel_CP_1635_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1635_elements(54);
      loadKernelChannel_CP_1635_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1635_elements(55);
      loadKernelChannel_CP_1635_elements(48) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1635_elements(49);
      loadKernelChannel_CP_1635_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1635_elements(58);
      loadKernelChannel_CP_1635_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1635_elements(59);
      loadKernelChannel_CP_1635_elements(50) <= phi_mux_reqs(1);
      phi_stmt_585_phi_seq_1885 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_585_phi_seq_1885") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1635_elements(43), 
          phi_sample_ack => loadKernelChannel_CP_1635_elements(44), 
          phi_update_req => loadKernelChannel_CP_1635_elements(45), 
          phi_update_ack => loadKernelChannel_CP_1635_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_1635_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1773_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_1635_elements(16);
        preds(1)  <= loadKernelChannel_CP_1635_elements(17);
        entry_tmerge_1773 : transition_merge -- 
          generic map(name => " entry_tmerge_1773")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_594_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_643_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_607_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_652_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_652_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_652_wire : std_logic_vector(63 downto 0);
    signal NOT_u1_u1_617_wire : std_logic_vector(0 downto 0);
    signal R_sh_start_541_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_541_scaled : std_logic_vector(13 downto 0);
    signal SHL_u16_u16_530_wire : std_logic_vector(15 downto 0);
    signal SHL_u16_u16_559_wire : std_logic_vector(15 downto 0);
    signal SUB_u64_u64_595_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_680_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_620_wire : std_logic_vector(0 downto 0);
    signal ULT_u64_u1_681_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_542_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_542_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_542_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_542_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_542_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_542_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_root_address : std_logic_vector(13 downto 0);
    signal ea1_554 : std_logic_vector(63 downto 0);
    signal ea2_562 : std_logic_vector(63 downto 0);
    signal ea3_568 : std_logic_vector(63 downto 0);
    signal fetch_addr_544 : std_logic_vector(31 downto 0);
    signal fetch_addr_655 : std_logic_vector(31 downto 0);
    signal fetch_val_585 : std_logic_vector(63 downto 0);
    signal fetch_val_616_delayed_13_0_669 : std_logic_vector(63 downto 0);
    signal first_fill_573 : std_logic_vector(0 downto 0);
    signal fn_608_delayed_7_0_658 : std_logic_vector(0 downto 0);
    signal fn_614_delayed_13_0_666 : std_logic_vector(0 downto 0);
    signal fn_646 : std_logic_vector(0 downto 0);
    signal fv_663 : std_logic_vector(63 downto 0);
    signal konst_529_wire_constant : std_logic_vector(15 downto 0);
    signal konst_535_wire_constant : std_logic_vector(63 downto 0);
    signal konst_558_wire_constant : std_logic_vector(15 downto 0);
    signal konst_571_wire_constant : std_logic_vector(63 downto 0);
    signal konst_591_wire_constant : std_logic_vector(63 downto 0);
    signal konst_593_wire_constant : std_logic_vector(63 downto 0);
    signal konst_596_wire_constant : std_logic_vector(63 downto 0);
    signal konst_601_wire_constant : std_logic_vector(63 downto 0);
    signal konst_642_wire_constant : std_logic_vector(63 downto 0);
    signal konst_644_wire_constant : std_logic_vector(63 downto 0);
    signal konst_651_wire_constant : std_logic_vector(63 downto 0);
    signal konst_679_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_548 : std_logic_vector(63 downto 0);
    signal my_fetch_548_588_buffered : std_logic_vector(63 downto 0);
    signal my_num1_598 : std_logic_vector(63 downto 0);
    signal mycount_581 : std_logic_vector(63 downto 0);
    signal nfetch_val_675 : std_logic_vector(63 downto 0);
    signal nfetch_val_675_587_buffered : std_logic_vector(63 downto 0);
    signal nmycount_603 : std_logic_vector(63 downto 0);
    signal nmycount_603_584_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_547_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_547_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_547_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_547_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_547_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_662_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_662_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_662_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_662_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_662_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_size_532 : std_logic_vector(15 downto 0);
    signal send_to_1_614 : std_logic_vector(0 downto 0);
    signal send_to_2_622 : std_logic_vector(0 downto 0);
    signal send_to_3_627 : std_logic_vector(0 downto 0);
    signal sh_start_537 : std_logic_vector(63 downto 0);
    signal start_add_583_buffered : std_logic_vector(63 downto 0);
    signal start_next_577 : std_logic_vector(7 downto 0);
    signal type_cast_552_wire : std_logic_vector(63 downto 0);
    signal type_cast_560_wire : std_logic_vector(63 downto 0);
    signal type_cast_566_wire : std_logic_vector(63 downto 0);
    signal var_val_609 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_542_constant_part_of_offset <= "00000000000000";
    array_obj_ref_542_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_542_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_542_resized_base_address <= "00000000000000";
    array_obj_ref_653_constant_part_of_offset <= "00000000000000";
    array_obj_ref_653_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_653_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_653_resized_base_address <= "00000000000000";
    konst_529_wire_constant <= "0000000000000001";
    konst_535_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_558_wire_constant <= "0000000000000001";
    konst_571_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_591_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_593_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_596_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_601_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_642_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    konst_644_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_651_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_679_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_547_word_offset_0 <= "00000000000000";
    ptr_deref_662_word_offset_0 <= "00000000000000";
    phi_stmt_581: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= start_add_583_buffered & nmycount_603_584_buffered;
      req <= phi_stmt_581_req_0 & phi_stmt_581_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_581",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_581_ack_0,
          idata => idata,
          odata => mycount_581,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_581
    phi_stmt_585: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nfetch_val_675_587_buffered & my_fetch_548_588_buffered;
      req <= phi_stmt_585_req_0 & phi_stmt_585_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_585",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_585_ack_0,
          idata => idata,
          odata => fetch_val_585,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_585
    -- flow-through select operator MUX_674_inst
    nfetch_val_675 <= fv_663 when (fn_614_delayed_13_0_666(0) /=  '0') else fetch_val_616_delayed_13_0_669;
    W_fetch_val_616_delayed_13_0_667_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_616_delayed_13_0_667_inst_req_0;
      W_fetch_val_616_delayed_13_0_667_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_616_delayed_13_0_667_inst_req_1;
      W_fetch_val_616_delayed_13_0_667_inst_ack_1<= rack(0);
      W_fetch_val_616_delayed_13_0_667_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_616_delayed_13_0_667_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_585,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_616_delayed_13_0_669,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_608_delayed_7_0_656_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_608_delayed_7_0_656_inst_req_0;
      W_fn_608_delayed_7_0_656_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_608_delayed_7_0_656_inst_req_1;
      W_fn_608_delayed_7_0_656_inst_ack_1<= rack(0);
      W_fn_608_delayed_7_0_656_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_608_delayed_7_0_656_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_608_delayed_7_0_658,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_614_delayed_13_0_664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_614_delayed_13_0_664_inst_req_0;
      W_fn_614_delayed_13_0_664_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_614_delayed_13_0_664_inst_req_1;
      W_fn_614_delayed_13_0_664_inst_ack_1<= rack(0);
      W_fn_614_delayed_13_0_664_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_614_delayed_13_0_664_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_614_delayed_13_0_666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_543_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_543_final_reg_req_0;
      addr_of_543_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_543_final_reg_req_1;
      addr_of_543_final_reg_ack_1<= rack(0);
      addr_of_543_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_543_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_542_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_544,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_654_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_654_final_reg_req_0;
      addr_of_654_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_654_final_reg_req_1;
      addr_of_654_final_reg_ack_1<= rack(0);
      addr_of_654_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_654_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_653_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_655,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_548_588_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_548_588_buf_req_0;
      my_fetch_548_588_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_548_588_buf_req_1;
      my_fetch_548_588_buf_ack_1<= rack(0);
      my_fetch_548_588_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_548_588_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_548_588_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_675_587_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_675_587_buf_req_0;
      nfetch_val_675_587_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_675_587_buf_req_1;
      nfetch_val_675_587_buf_ack_1<= rack(0);
      nfetch_val_675_587_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_675_587_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_675,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_675_587_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_603_584_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_603_584_buf_req_0;
      nmycount_603_584_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_603_584_buf_req_1;
      nmycount_603_584_buf_ack_1<= rack(0);
      nmycount_603_584_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_603_584_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_603,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_603_584_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_583_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_583_buf_req_0;
      start_add_583_buf_ack_0<= wack(0);
      rreq(0) <= start_add_583_buf_req_1;
      start_add_583_buf_ack_1<= rack(0);
      start_add_583_buf : InterlockBuffer generic map ( -- 
        name => "start_add_583_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_583_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_552_inst
    process(row_size_532) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_532(15 downto 0);
      type_cast_552_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_560_inst
    process(SHL_u16_u16_559_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := SHL_u16_u16_559_wire(15 downto 0);
      type_cast_560_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_566_inst
    process(row_size_532) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_532(15 downto 0);
      type_cast_566_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_608_inst
    process(LSHR_u64_u64_607_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := LSHR_u64_u64_607_wire(7 downto 0);
      var_val_609 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_542_index_1_rename
    process(R_sh_start_541_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_541_resized;
      ov(13 downto 0) := iv;
      R_sh_start_541_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_542_index_1_resize
    process(sh_start_537) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_537;
      ov := iv(13 downto 0);
      R_sh_start_541_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_542_root_address_inst
    process(array_obj_ref_542_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_542_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_542_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_653_index_1_rename
    process(LSHR_u64_u64_652_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_652_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_652_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_653_index_1_resize
    process(LSHR_u64_u64_652_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_652_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_652_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_653_root_address_inst
    process(array_obj_ref_653_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_653_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_653_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_547_addr_0
    process(ptr_deref_547_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_547_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_547_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_547_base_resize
    process(fetch_addr_544) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_544;
      ov := iv(13 downto 0);
      ptr_deref_547_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_547_gather_scatter
    process(ptr_deref_547_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_547_data_0;
      ov(63 downto 0) := iv;
      my_fetch_548 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_547_root_address_inst
    process(ptr_deref_547_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_547_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_547_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_662_addr_0
    process(ptr_deref_662_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_662_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_662_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_662_base_resize
    process(fetch_addr_655) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_655;
      ov := iv(13 downto 0);
      ptr_deref_662_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_662_gather_scatter
    process(ptr_deref_662_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_662_data_0;
      ov(63 downto 0) := iv;
      fv_663 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_662_root_address_inst
    process(ptr_deref_662_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_662_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_662_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_579_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_681_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_579_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_579_branch_req_0,
          ack0 => do_while_stmt_579_branch_ack_0,
          ack1 => do_while_stmt_579_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_531_inst
    process(num_chl_buffer, SHL_u16_u16_530_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_chl_buffer, SHL_u16_u16_530_wire, tmp_var);
      row_size_532 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_553_inst
    process(start_add_buffer, type_cast_552_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_552_wire, tmp_var);
      ea1_554 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_561_inst
    process(start_add_buffer, type_cast_560_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_560_wire, tmp_var);
      ea2_562 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_567_inst
    process(ea2_562, type_cast_566_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ea2_562, type_cast_566_wire, tmp_var);
      ea3_568 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_602_inst
    process(mycount_581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_581, konst_601_wire_constant, tmp_var);
      nmycount_603 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_621_inst
    process(NOT_u1_u1_617_wire, ULT_u64_u1_620_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_617_wire, ULT_u64_u1_620_wire, tmp_var);
      send_to_2_622 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_594_inst
    process(mycount_581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_581, konst_593_wire_constant, tmp_var);
      AND_u64_u64_594_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_643_inst
    process(nmycount_603) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_603, konst_642_wire_constant, tmp_var);
      AND_u64_u64_643_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_572_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_571_wire_constant, tmp_var);
      first_fill_573 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_645_inst
    process(AND_u64_u64_643_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_643_wire, konst_644_wire_constant, tmp_var);
      fn_646 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_536_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_535_wire_constant, tmp_var);
      sh_start_537 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_607_inst
    process(fetch_val_585, my_num1_598) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_585, my_num1_598, tmp_var);
      LSHR_u64_u64_607_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_652_inst
    process(nmycount_603) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_603, konst_651_wire_constant, tmp_var);
      LSHR_u64_u64_652_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_617_inst
    process(send_to_1_614) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", send_to_1_614, tmp_var);
      NOT_u1_u1_617_wire <= tmp_var; -- 
    end process;
    -- binary operator SHL_u16_u16_530_inst
    process(num_chl_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(num_chl_buffer, konst_529_wire_constant, tmp_var);
      SHL_u16_u16_530_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_559_inst
    process(row_size_532) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(row_size_532, konst_558_wire_constant, tmp_var);
      SHL_u16_u16_559_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_597_inst
    process(SUB_u64_u64_595_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_595_wire, konst_596_wire_constant, tmp_var);
      my_num1_598 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_595_inst
    process(konst_591_wire_constant, AND_u64_u64_594_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_591_wire_constant, AND_u64_u64_594_wire, tmp_var);
      SUB_u64_u64_595_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_680_inst
    process(ea3_568) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(ea3_568, konst_679_wire_constant, tmp_var);
      SUB_u64_u64_680_wire <= tmp_var; --
    end process;
    -- binary operator UGE_u64_u1_626_inst
    process(mycount_581, ea2_562) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(mycount_581, ea2_562, tmp_var);
      send_to_3_627 <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_613_inst
    process(mycount_581, ea1_554) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_581, ea1_554, tmp_var);
      send_to_1_614 <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_620_inst
    process(mycount_581, ea2_562) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_581, ea2_562, tmp_var);
      ULT_u64_u1_620_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_681_inst
    process(mycount_581, SUB_u64_u64_680_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_581, SUB_u64_u64_680_wire, tmp_var);
      ULT_u64_u1_681_wire <= tmp_var; --
    end process;
    -- shared split operator group (23) : array_obj_ref_542_index_offset 
    ApIntAdd_group_23: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_541_scaled;
      array_obj_ref_542_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_542_index_offset_req_0;
      array_obj_ref_542_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_542_index_offset_req_1;
      array_obj_ref_542_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_23_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : array_obj_ref_653_index_offset 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_652_scaled;
      array_obj_ref_653_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_653_index_offset_req_0;
      array_obj_ref_653_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_653_index_offset_req_1;
      array_obj_ref_653_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_24_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared load operator group (0) : ptr_deref_547_load_0 ptr_deref_662_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_547_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_662_load_0_req_0;
      ptr_deref_547_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_662_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_547_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_662_load_0_req_1;
      ptr_deref_547_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_662_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_608_delayed_7_0_658(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_547_word_address_0 & ptr_deref_662_word_address_0;
      ptr_deref_547_data_0 <= data_out(127 downto 64);
      ptr_deref_662_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_576_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_576_inst_req_0;
      RPIPE_input_done_pipe_576_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_576_inst_req_1;
      RPIPE_input_done_pipe_576_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_573(0);
      start_next_577 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_629_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_629_inst_req_0;
      WPIPE_kernel_pipe1_629_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_629_inst_req_1;
      WPIPE_kernel_pipe1_629_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_614(0);
      data_in <= var_val_609;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe2_633_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe2_633_inst_req_0;
      WPIPE_kernel_pipe2_633_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe2_633_inst_req_1;
      WPIPE_kernel_pipe2_633_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_622(0);
      data_in <= var_val_609;
      kernel_pipe2_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe2", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe2_pipe_write_req(0),
          oack => kernel_pipe2_pipe_write_ack(0),
          odata => kernel_pipe2_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_kernel_pipe3_637_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe3_637_inst_req_0;
      WPIPE_kernel_pipe3_637_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe3_637_inst_req_1;
      WPIPE_kernel_pipe3_637_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_627(0);
      data_in <= var_val_609;
      kernel_pipe3_write_2_gI: SplitGuardInterface generic map(name => "kernel_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "kernel_pipe3", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe3_pipe_write_req(0),
          oack => kernel_pipe3_pipe_write_ack(0),
          odata => kernel_pipe3_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_size_pipe_683_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_683_inst_req_0;
      WPIPE_size_pipe_683_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_683_inst_req_1;
      WPIPE_size_pipe_683_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= num_chl_buffer;
      size_pipe_write_3_gI: SplitGuardInterface generic map(name => "size_pipe_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_3: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendB is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendB;
architecture sendB_arch of sendB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendB_CP_2093_start: Boolean;
  signal sendB_CP_2093_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_1095_branch_req_0 : boolean;
  signal ptr_deref_981_store_0_ack_0 : boolean;
  signal if_stmt_702_branch_req_0 : boolean;
  signal type_cast_992_inst_req_0 : boolean;
  signal type_cast_742_inst_ack_0 : boolean;
  signal if_stmt_702_branch_ack_1 : boolean;
  signal type_cast_742_inst_req_0 : boolean;
  signal type_cast_742_inst_req_1 : boolean;
  signal ptr_deref_981_store_0_req_0 : boolean;
  signal type_cast_742_inst_ack_1 : boolean;
  signal if_stmt_702_branch_ack_0 : boolean;
  signal ptr_deref_1065_store_0_ack_0 : boolean;
  signal type_cast_992_inst_ack_0 : boolean;
  signal type_cast_992_inst_req_1 : boolean;
  signal array_obj_ref_1179_final_reg_req_0 : boolean;
  signal ptr_deref_1086_store_0_ack_0 : boolean;
  signal type_cast_992_inst_ack_1 : boolean;
  signal if_stmt_1095_branch_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1137_inst_req_0 : boolean;
  signal array_obj_ref_1179_index_offset_ack_0 : boolean;
  signal if_stmt_1095_branch_ack_0 : boolean;
  signal array_obj_ref_1179_final_reg_req_1 : boolean;
  signal array_obj_ref_1179_final_reg_ack_1 : boolean;
  signal array_obj_ref_1179_final_reg_ack_0 : boolean;
  signal if_stmt_1146_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1137_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1137_inst_ack_0 : boolean;
  signal array_obj_ref_1179_index_offset_req_0 : boolean;
  signal type_cast_1034_inst_req_0 : boolean;
  signal if_stmt_1146_branch_ack_1 : boolean;
  signal ptr_deref_1002_store_0_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1137_inst_ack_1 : boolean;
  signal type_cast_1104_inst_req_1 : boolean;
  signal type_cast_1104_inst_ack_1 : boolean;
  signal ptr_deref_1086_store_0_req_1 : boolean;
  signal type_cast_1034_inst_ack_0 : boolean;
  signal if_stmt_1146_branch_req_0 : boolean;
  signal ptr_deref_981_store_0_req_1 : boolean;
  signal array_obj_ref_764_index_offset_req_0 : boolean;
  signal array_obj_ref_764_index_offset_ack_0 : boolean;
  signal array_obj_ref_764_index_offset_req_1 : boolean;
  signal array_obj_ref_764_index_offset_ack_1 : boolean;
  signal addr_of_765_final_reg_req_0 : boolean;
  signal addr_of_765_final_reg_ack_0 : boolean;
  signal addr_of_765_final_reg_req_1 : boolean;
  signal addr_of_765_final_reg_ack_1 : boolean;
  signal ptr_deref_769_load_0_req_0 : boolean;
  signal ptr_deref_769_load_0_ack_0 : boolean;
  signal ptr_deref_769_load_0_req_1 : boolean;
  signal ptr_deref_769_load_0_ack_1 : boolean;
  signal type_cast_773_inst_req_0 : boolean;
  signal type_cast_773_inst_ack_0 : boolean;
  signal type_cast_773_inst_req_1 : boolean;
  signal type_cast_773_inst_ack_1 : boolean;
  signal type_cast_783_inst_req_0 : boolean;
  signal type_cast_783_inst_ack_0 : boolean;
  signal type_cast_783_inst_req_1 : boolean;
  signal type_cast_783_inst_ack_1 : boolean;
  signal type_cast_793_inst_req_0 : boolean;
  signal type_cast_793_inst_ack_0 : boolean;
  signal type_cast_793_inst_req_1 : boolean;
  signal type_cast_793_inst_ack_1 : boolean;
  signal type_cast_803_inst_req_0 : boolean;
  signal type_cast_803_inst_ack_0 : boolean;
  signal type_cast_803_inst_req_1 : boolean;
  signal type_cast_803_inst_ack_1 : boolean;
  signal type_cast_813_inst_req_0 : boolean;
  signal type_cast_813_inst_ack_0 : boolean;
  signal type_cast_813_inst_req_1 : boolean;
  signal type_cast_813_inst_ack_1 : boolean;
  signal type_cast_823_inst_req_0 : boolean;
  signal type_cast_823_inst_ack_0 : boolean;
  signal type_cast_823_inst_req_1 : boolean;
  signal type_cast_823_inst_ack_1 : boolean;
  signal type_cast_833_inst_req_0 : boolean;
  signal type_cast_833_inst_ack_0 : boolean;
  signal type_cast_833_inst_req_1 : boolean;
  signal type_cast_833_inst_ack_1 : boolean;
  signal type_cast_843_inst_req_0 : boolean;
  signal type_cast_843_inst_ack_0 : boolean;
  signal type_cast_843_inst_req_1 : boolean;
  signal type_cast_843_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_845_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_845_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_845_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_845_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_848_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_848_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_848_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_848_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_851_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_851_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_851_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_851_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_854_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_854_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_854_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_854_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_857_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_857_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_857_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_857_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_860_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_860_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_860_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_860_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_863_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_863_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_863_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_863_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_866_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_866_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_866_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_866_inst_ack_1 : boolean;
  signal ptr_deref_1086_store_0_req_0 : boolean;
  signal type_cast_1013_inst_ack_1 : boolean;
  signal ptr_deref_1023_store_0_ack_1 : boolean;
  signal if_stmt_880_branch_req_0 : boolean;
  signal type_cast_1013_inst_req_1 : boolean;
  signal ptr_deref_1023_store_0_req_1 : boolean;
  signal if_stmt_880_branch_ack_1 : boolean;
  signal if_stmt_880_branch_ack_0 : boolean;
  signal ptr_deref_1065_store_0_req_0 : boolean;
  signal type_cast_896_inst_req_0 : boolean;
  signal type_cast_896_inst_ack_0 : boolean;
  signal type_cast_896_inst_req_1 : boolean;
  signal type_cast_896_inst_ack_1 : boolean;
  signal type_cast_1104_inst_ack_0 : boolean;
  signal type_cast_1076_inst_ack_1 : boolean;
  signal type_cast_1076_inst_req_1 : boolean;
  signal if_stmt_920_branch_req_0 : boolean;
  signal if_stmt_920_branch_ack_1 : boolean;
  signal if_stmt_920_branch_ack_0 : boolean;
  signal type_cast_929_inst_req_0 : boolean;
  signal type_cast_929_inst_ack_0 : boolean;
  signal type_cast_1076_inst_ack_0 : boolean;
  signal type_cast_929_inst_req_1 : boolean;
  signal type_cast_929_inst_ack_1 : boolean;
  signal type_cast_1104_inst_req_0 : boolean;
  signal type_cast_1055_inst_ack_1 : boolean;
  signal type_cast_1055_inst_req_1 : boolean;
  signal type_cast_1013_inst_ack_0 : boolean;
  signal type_cast_1013_inst_req_0 : boolean;
  signal ptr_deref_1023_store_0_ack_0 : boolean;
  signal array_obj_ref_935_index_offset_req_0 : boolean;
  signal array_obj_ref_935_index_offset_ack_0 : boolean;
  signal array_obj_ref_935_index_offset_req_1 : boolean;
  signal array_obj_ref_935_index_offset_ack_1 : boolean;
  signal type_cast_1076_inst_req_0 : boolean;
  signal addr_of_936_final_reg_req_0 : boolean;
  signal addr_of_936_final_reg_ack_0 : boolean;
  signal ptr_deref_1023_store_0_req_0 : boolean;
  signal addr_of_936_final_reg_req_1 : boolean;
  signal addr_of_936_final_reg_ack_1 : boolean;
  signal type_cast_1055_inst_ack_0 : boolean;
  signal type_cast_1055_inst_req_0 : boolean;
  signal ptr_deref_940_load_0_req_0 : boolean;
  signal ptr_deref_940_load_0_ack_0 : boolean;
  signal ptr_deref_940_load_0_req_1 : boolean;
  signal ptr_deref_940_load_0_ack_1 : boolean;
  signal ptr_deref_1002_store_0_ack_1 : boolean;
  signal array_obj_ref_1179_index_offset_ack_1 : boolean;
  signal ptr_deref_1044_store_0_ack_1 : boolean;
  signal ptr_deref_1002_store_0_req_1 : boolean;
  signal type_cast_950_inst_req_0 : boolean;
  signal type_cast_950_inst_ack_0 : boolean;
  signal type_cast_950_inst_req_1 : boolean;
  signal type_cast_950_inst_ack_1 : boolean;
  signal array_obj_ref_1179_index_offset_req_1 : boolean;
  signal ptr_deref_1044_store_0_req_1 : boolean;
  signal ptr_deref_1044_store_0_ack_0 : boolean;
  signal type_cast_1034_inst_ack_1 : boolean;
  signal ptr_deref_960_store_0_req_0 : boolean;
  signal ptr_deref_960_store_0_ack_0 : boolean;
  signal ptr_deref_1065_store_0_ack_1 : boolean;
  signal ptr_deref_960_store_0_req_1 : boolean;
  signal ptr_deref_960_store_0_ack_1 : boolean;
  signal ptr_deref_1086_store_0_ack_1 : boolean;
  signal ptr_deref_1044_store_0_req_0 : boolean;
  signal ptr_deref_1065_store_0_req_1 : boolean;
  signal ptr_deref_1002_store_0_ack_0 : boolean;
  signal type_cast_971_inst_req_0 : boolean;
  signal type_cast_1034_inst_req_1 : boolean;
  signal type_cast_971_inst_ack_0 : boolean;
  signal type_cast_971_inst_req_1 : boolean;
  signal type_cast_971_inst_ack_1 : boolean;
  signal ptr_deref_981_store_0_ack_1 : boolean;
  signal ptr_deref_1183_load_0_req_0 : boolean;
  signal ptr_deref_1183_load_0_ack_0 : boolean;
  signal ptr_deref_1183_load_0_req_1 : boolean;
  signal ptr_deref_1183_load_0_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1185_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1185_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1185_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1185_inst_ack_1 : boolean;
  signal if_stmt_1193_branch_req_0 : boolean;
  signal if_stmt_1193_branch_ack_1 : boolean;
  signal if_stmt_1193_branch_ack_0 : boolean;
  signal phi_stmt_752_req_0 : boolean;
  signal type_cast_758_inst_req_0 : boolean;
  signal type_cast_758_inst_ack_0 : boolean;
  signal type_cast_758_inst_req_1 : boolean;
  signal type_cast_758_inst_ack_1 : boolean;
  signal phi_stmt_752_req_1 : boolean;
  signal phi_stmt_752_ack_0 : boolean;
  signal phi_stmt_900_req_1 : boolean;
  signal type_cast_903_inst_req_0 : boolean;
  signal type_cast_903_inst_ack_0 : boolean;
  signal type_cast_903_inst_req_1 : boolean;
  signal type_cast_903_inst_ack_1 : boolean;
  signal phi_stmt_900_req_0 : boolean;
  signal phi_stmt_900_ack_0 : boolean;
  signal phi_stmt_1161_req_1 : boolean;
  signal type_cast_1164_inst_req_0 : boolean;
  signal type_cast_1164_inst_ack_0 : boolean;
  signal type_cast_1164_inst_req_1 : boolean;
  signal type_cast_1164_inst_ack_1 : boolean;
  signal phi_stmt_1161_req_0 : boolean;
  signal phi_stmt_1161_ack_0 : boolean;
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(2 downto 0);
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendB_CP_2093_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2093_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendB_CP_2093_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2093_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendB_CP_2093: Block -- control-path 
    signal sendB_CP_2093_elements: BooleanArray(145 downto 0);
    -- 
  begin -- 
    sendB_CP_2093_elements(0) <= sendB_CP_2093_start;
    sendB_CP_2093_symbol <= sendB_CP_2093_elements(145);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 branch_block_stmt_689/assign_stmt_695_to_assign_stmt_701/$exit
      -- CP-element group 0: 	 branch_block_stmt_689/assign_stmt_695_to_assign_stmt_701/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_else_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_689/R_cmp76_703_place
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_689/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/branch_block_stmt_689__entry__
      -- CP-element group 0: 	 branch_block_stmt_689/assign_stmt_695_to_assign_stmt_701__entry__
      -- CP-element group 0: 	 branch_block_stmt_689/assign_stmt_695_to_assign_stmt_701__exit__
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702__entry__
      -- 
    branch_req_2167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(0), ack => if_stmt_702_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	3 
    -- CP-element group 1: 	4 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_689/if_stmt_702_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_689/if_stmt_702_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_689/entry_bbx_xnph78
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/$entry
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_update_start_
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_689/merge_stmt_708__exit__
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749__entry__
      -- CP-element group 1: 	 branch_block_stmt_689/entry_bbx_xnph78_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_689/entry_bbx_xnph78_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_689/merge_stmt_708_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_689/merge_stmt_708_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_689/merge_stmt_708_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_689/merge_stmt_708_PhiAck/dummy
      -- 
    if_choice_transition_2172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_702_branch_ack_1, ack => sendB_CP_2093_elements(1)); -- 
    rr_2189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(1), ack => type_cast_742_inst_req_0); -- 
    cr_2194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(1), ack => type_cast_742_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	133 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_689/if_stmt_702_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_689/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_689/if_stmt_702_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_900/$entry
      -- CP-element group 2: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/$entry
      -- 
    else_choice_transition_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_702_branch_ack_0, ack => sendB_CP_2093_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_sample_completed_
      -- 
    ra_2190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_742_inst_ack_0, ack => sendB_CP_2093_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	127 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_689/bbx_xnph78_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/$exit
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749/type_cast_742_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_749__exit__
      -- CP-element group 4: 	 branch_block_stmt_689/bbx_xnph78_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_689/bbx_xnph78_forx_xbody_PhiReq/phi_stmt_752/$entry
      -- CP-element group 4: 	 branch_block_stmt_689/bbx_xnph78_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/$entry
      -- 
    ca_2195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_742_inst_ack_1, ack => sendB_CP_2093_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	132 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_final_index_sum_regn_Sample/ack
      -- 
    ack_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_764_index_offset_ack_0, ack => sendB_CP_2093_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	132 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_request/req
      -- 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_764_index_offset_ack_1, ack => sendB_CP_2093_elements(6)); -- 
    req_2238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(6), ack => addr_of_765_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_request/$exit
      -- CP-element group 7: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_request/ack
      -- 
    ack_2239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_765_final_reg_ack_0, ack => sendB_CP_2093_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	132 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Sample/word_access_start/word_0/rr
      -- 
    ack_2244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_765_final_reg_ack_1, ack => sendB_CP_2093_elements(8)); -- 
    rr_2277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(8), ack => ptr_deref_769_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Sample/word_access_start/word_0/ra
      -- 
    ra_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_769_load_0_ack_0, ack => sendB_CP_2093_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	132 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	21 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	25 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/ptr_deref_769_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/ptr_deref_769_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/ptr_deref_769_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/ptr_deref_769_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_Sample/rr
      -- 
    ca_2289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_769_load_0_ack_1, ack => sendB_CP_2093_elements(10)); -- 
    rr_2302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(10), ack => type_cast_773_inst_req_0); -- 
    rr_2316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(10), ack => type_cast_783_inst_req_0); -- 
    rr_2330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(10), ack => type_cast_793_inst_req_0); -- 
    rr_2344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(10), ack => type_cast_803_inst_req_0); -- 
    rr_2358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(10), ack => type_cast_813_inst_req_0); -- 
    rr_2372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(10), ack => type_cast_823_inst_req_0); -- 
    rr_2386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(10), ack => type_cast_833_inst_req_0); -- 
    rr_2400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(10), ack => type_cast_843_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_Sample/ra
      -- 
    ra_2303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_773_inst_ack_0, ack => sendB_CP_2093_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	132 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	47 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_Update/ca
      -- 
    ca_2308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_773_inst_ack_1, ack => sendB_CP_2093_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_Sample/ra
      -- 
    ra_2317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_783_inst_ack_0, ack => sendB_CP_2093_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	132 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	44 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_Update/ca
      -- 
    ca_2322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_783_inst_ack_1, ack => sendB_CP_2093_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_Sample/ra
      -- 
    ra_2331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_0, ack => sendB_CP_2093_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	132 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_Update/ca
      -- 
    ca_2336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_1, ack => sendB_CP_2093_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_Sample/ra
      -- 
    ra_2345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_803_inst_ack_0, ack => sendB_CP_2093_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	132 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	38 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_Update/ca
      -- 
    ca_2350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_803_inst_ack_1, ack => sendB_CP_2093_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_Sample/ra
      -- 
    ra_2359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_813_inst_ack_0, ack => sendB_CP_2093_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	132 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	35 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_Update/ca
      -- 
    ca_2364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_813_inst_ack_1, ack => sendB_CP_2093_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	10 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_Sample/ra
      -- 
    ra_2373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_823_inst_ack_0, ack => sendB_CP_2093_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	132 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	32 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_Update/ca
      -- 
    ca_2378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_823_inst_ack_1, ack => sendB_CP_2093_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_Sample/ra
      -- 
    ra_2387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_0, ack => sendB_CP_2093_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	132 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_Update/ca
      -- 
    ca_2392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_1, ack => sendB_CP_2093_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_Sample/ra
      -- 
    ra_2401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_0, ack => sendB_CP_2093_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	132 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_Sample/req
      -- 
    ca_2406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_1, ack => sendB_CP_2093_elements(26)); -- 
    req_2414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(26), ack => WPIPE_maxpool_output_pipe_845_inst_req_0); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_update_start_
      -- CP-element group 27: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_Update/req
      -- 
    ack_2415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_845_inst_ack_0, ack => sendB_CP_2093_elements(27)); -- 
    req_2419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(27), ack => WPIPE_maxpool_output_pipe_845_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_845_Update/ack
      -- 
    ack_2420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_845_inst_ack_1, ack => sendB_CP_2093_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_Sample/req
      -- 
    req_2428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(29), ack => WPIPE_maxpool_output_pipe_848_inst_req_0); -- 
    sendB_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(24) & sendB_CP_2093_elements(28);
      gj_sendB_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_update_start_
      -- CP-element group 30: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_Update/req
      -- 
    ack_2429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_848_inst_ack_0, ack => sendB_CP_2093_elements(30)); -- 
    req_2433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(30), ack => WPIPE_maxpool_output_pipe_848_inst_req_1); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_848_Update/ack
      -- 
    ack_2434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_848_inst_ack_1, ack => sendB_CP_2093_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	22 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_Sample/req
      -- 
    req_2442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(32), ack => WPIPE_maxpool_output_pipe_851_inst_req_0); -- 
    sendB_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(22) & sendB_CP_2093_elements(31);
      gj_sendB_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_update_start_
      -- CP-element group 33: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_Update/req
      -- 
    ack_2443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_851_inst_ack_0, ack => sendB_CP_2093_elements(33)); -- 
    req_2447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(33), ack => WPIPE_maxpool_output_pipe_851_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_851_Update/ack
      -- 
    ack_2448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_851_inst_ack_1, ack => sendB_CP_2093_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	20 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_Sample/req
      -- 
    req_2456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(35), ack => WPIPE_maxpool_output_pipe_854_inst_req_0); -- 
    sendB_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(20) & sendB_CP_2093_elements(34);
      gj_sendB_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_update_start_
      -- CP-element group 36: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_Update/req
      -- 
    ack_2457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_854_inst_ack_0, ack => sendB_CP_2093_elements(36)); -- 
    req_2461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(36), ack => WPIPE_maxpool_output_pipe_854_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_854_Update/ack
      -- 
    ack_2462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_854_inst_ack_1, ack => sendB_CP_2093_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	18 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_Sample/req
      -- 
    req_2470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(38), ack => WPIPE_maxpool_output_pipe_857_inst_req_0); -- 
    sendB_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(18) & sendB_CP_2093_elements(37);
      gj_sendB_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_update_start_
      -- CP-element group 39: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_Update/req
      -- 
    ack_2471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_857_inst_ack_0, ack => sendB_CP_2093_elements(39)); -- 
    req_2475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(39), ack => WPIPE_maxpool_output_pipe_857_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_857_Update/ack
      -- 
    ack_2476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_857_inst_ack_1, ack => sendB_CP_2093_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_Sample/req
      -- 
    req_2484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(41), ack => WPIPE_maxpool_output_pipe_860_inst_req_0); -- 
    sendB_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(16) & sendB_CP_2093_elements(40);
      gj_sendB_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_update_start_
      -- CP-element group 42: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_Update/req
      -- 
    ack_2485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_860_inst_ack_0, ack => sendB_CP_2093_elements(42)); -- 
    req_2489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(42), ack => WPIPE_maxpool_output_pipe_860_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_860_Update/ack
      -- 
    ack_2490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_860_inst_ack_1, ack => sendB_CP_2093_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	14 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_Sample/req
      -- 
    req_2498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(44), ack => WPIPE_maxpool_output_pipe_863_inst_req_0); -- 
    sendB_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(14) & sendB_CP_2093_elements(43);
      gj_sendB_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_update_start_
      -- CP-element group 45: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_Update/req
      -- 
    ack_2499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_863_inst_ack_0, ack => sendB_CP_2093_elements(45)); -- 
    req_2503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(45), ack => WPIPE_maxpool_output_pipe_863_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_863_Update/ack
      -- 
    ack_2504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_863_inst_ack_1, ack => sendB_CP_2093_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	12 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_Sample/req
      -- 
    req_2512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(47), ack => WPIPE_maxpool_output_pipe_866_inst_req_0); -- 
    sendB_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(12) & sendB_CP_2093_elements(46);
      gj_sendB_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_update_start_
      -- CP-element group 48: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_Update/req
      -- 
    ack_2513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_866_inst_ack_0, ack => sendB_CP_2093_elements(48)); -- 
    req_2517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(48), ack => WPIPE_maxpool_output_pipe_866_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/WPIPE_maxpool_output_pipe_866_Update/ack
      -- 
    ack_2518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_866_inst_ack_1, ack => sendB_CP_2093_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_689/if_stmt_880__entry__
      -- CP-element group 50: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879__exit__
      -- CP-element group 50: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/$exit
      -- CP-element group 50: 	 branch_block_stmt_689/if_stmt_880_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_689/if_stmt_880_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_689/if_stmt_880_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_689/if_stmt_880_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_689/R_exitcond_881_place
      -- CP-element group 50: 	 branch_block_stmt_689/if_stmt_880_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_689/if_stmt_880_else_link/$entry
      -- 
    branch_req_2526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(50), ack => if_stmt_880_branch_req_0); -- 
    sendB_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(5) & sendB_CP_2093_elements(49);
      gj_sendB_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: 	54 
    -- CP-element group 51:  members (18) 
      -- CP-element group 51: 	 branch_block_stmt_689/merge_stmt_886__exit__
      -- CP-element group 51: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897__entry__
      -- CP-element group 51: 	 branch_block_stmt_689/if_stmt_880_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_689/if_stmt_880_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_689/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 51: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/$entry
      -- CP-element group 51: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_update_start_
      -- CP-element group 51: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_689/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_689/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_689/merge_stmt_886_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_689/merge_stmt_886_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_689/merge_stmt_886_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_689/merge_stmt_886_PhiAck/dummy
      -- 
    if_choice_transition_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_880_branch_ack_1, ack => sendB_CP_2093_elements(51)); -- 
    rr_2548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(51), ack => type_cast_896_inst_req_0); -- 
    cr_2553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(51), ack => type_cast_896_inst_req_1); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	128 
    -- CP-element group 52: 	129 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_689/if_stmt_880_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/if_stmt_880_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_880_branch_ack_0, ack => sendB_CP_2093_elements(52)); -- 
    rr_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => type_cast_758_inst_req_0); -- 
    cr_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => type_cast_758_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_Sample/ra
      -- 
    ra_2549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_896_inst_ack_0, ack => sendB_CP_2093_elements(53)); -- 
    -- CP-element group 54:  fork  transition  place  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	134 
    -- CP-element group 54: 	135 
    -- CP-element group 54:  members (15) 
      -- CP-element group 54: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 54: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897__exit__
      -- CP-element group 54: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/$exit
      -- CP-element group 54: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_689/assign_stmt_893_to_assign_stmt_897/type_cast_896_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/$entry
      -- CP-element group 54: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/$entry
      -- CP-element group 54: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/$entry
      -- CP-element group 54: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/SplitProtocol/$entry
      -- CP-element group 54: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/SplitProtocol/Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/SplitProtocol/Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/SplitProtocol/Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/SplitProtocol/Update/cr
      -- 
    ca_2554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_896_inst_ack_1, ack => sendB_CP_2093_elements(54)); -- 
    rr_3447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(54), ack => type_cast_903_inst_req_0); -- 
    cr_3452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(54), ack => type_cast_903_inst_req_1); -- 
    -- CP-element group 55:  transition  place  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	138 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	145 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_689/if_stmt_920_if_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_689/if_stmt_920_if_link/if_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_689/forx_xend_sendRemainingElementsx_xexit
      -- CP-element group 55: 	 branch_block_stmt_689/forx_xend_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_689/forx_xend_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_920_branch_ack_1, ack => sendB_CP_2093_elements(55)); -- 
    -- CP-element group 56:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	138 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56: 	59 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	62 
    -- CP-element group 56: 	64 
    -- CP-element group 56: 	66 
    -- CP-element group 56: 	67 
    -- CP-element group 56: 	69 
    -- CP-element group 56: 	71 
    -- CP-element group 56: 	72 
    -- CP-element group 56: 	74 
    -- CP-element group 56: 	76 
    -- CP-element group 56: 	77 
    -- CP-element group 56: 	79 
    -- CP-element group 56: 	81 
    -- CP-element group 56: 	82 
    -- CP-element group 56: 	84 
    -- CP-element group 56: 	86 
    -- CP-element group 56: 	87 
    -- CP-element group 56: 	89 
    -- CP-element group 56: 	91 
    -- CP-element group 56: 	92 
    -- CP-element group 56: 	94 
    -- CP-element group 56: 	96 
    -- CP-element group 56: 	97 
    -- CP-element group 56: 	99 
    -- CP-element group 56:  members (210) 
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094__entry__
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_689/merge_stmt_926__exit__
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/if_stmt_920_else_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_689/if_stmt_920_else_link/else_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_689/forx_xend_ifx_xthen
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_final_index_sum_regn_update_start
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_final_index_sum_regn_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_final_index_sum_regn_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_final_index_sum_regn_Update/req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_complete/req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_update_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_689/forx_xend_ifx_xthen_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/forx_xend_ifx_xthen_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/merge_stmt_926_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_689/merge_stmt_926_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/merge_stmt_926_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/merge_stmt_926_PhiAck/dummy
      -- 
    else_choice_transition_2574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_920_branch_ack_0, ack => sendB_CP_2093_elements(56)); -- 
    cr_2830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => type_cast_992_inst_req_1); -- 
    cr_3136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => ptr_deref_1086_store_0_req_1); -- 
    cr_2816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => ptr_deref_981_store_0_req_1); -- 
    cr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => type_cast_1013_inst_req_1); -- 
    cr_2944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => ptr_deref_1023_store_0_req_1); -- 
    cr_3086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => type_cast_1076_inst_req_1); -- 
    rr_2587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => type_cast_929_inst_req_0); -- 
    cr_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => type_cast_929_inst_req_1); -- 
    cr_3022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => type_cast_1055_inst_req_1); -- 
    req_2618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => array_obj_ref_935_index_offset_req_0); -- 
    req_2623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => array_obj_ref_935_index_offset_req_1); -- 
    req_2638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => addr_of_936_final_reg_req_1); -- 
    cr_2683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => ptr_deref_940_load_0_req_1); -- 
    cr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => ptr_deref_1002_store_0_req_1); -- 
    cr_2702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => type_cast_950_inst_req_1); -- 
    cr_3008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => ptr_deref_1044_store_0_req_1); -- 
    cr_2752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => ptr_deref_960_store_0_req_1); -- 
    cr_3072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => ptr_deref_1065_store_0_req_1); -- 
    cr_2958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => type_cast_1034_inst_req_1); -- 
    cr_2766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => type_cast_971_inst_req_1); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_Sample/ra
      -- 
    ra_2588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_929_inst_ack_0, ack => sendB_CP_2093_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	106 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_929_Update/ca
      -- 
    ca_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_929_inst_ack_1, ack => sendB_CP_2093_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	56 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	106 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_final_index_sum_regn_Sample/ack
      -- 
    ack_2619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_935_index_offset_ack_0, ack => sendB_CP_2093_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/array_obj_ref_935_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_request/req
      -- 
    ack_2624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_935_index_offset_ack_1, ack => sendB_CP_2093_elements(60)); -- 
    req_2633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(60), ack => addr_of_936_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_request/ack
      -- 
    ack_2634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_936_final_reg_ack_0, ack => sendB_CP_2093_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	56 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (24) 
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/addr_of_936_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_word_addrgen/root_register_ack
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Sample/word_access_start/$entry
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Sample/word_access_start/word_0/$entry
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Sample/word_access_start/word_0/rr
      -- 
    ack_2639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_936_final_reg_ack_1, ack => sendB_CP_2093_elements(62)); -- 
    rr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(62), ack => ptr_deref_940_load_0_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Sample/word_access_start/$exit
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Sample/word_access_start/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Sample/word_access_start/word_0/ra
      -- 
    ra_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_940_load_0_ack_0, ack => sendB_CP_2093_elements(63)); -- 
    -- CP-element group 64:  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	56 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	70 
    -- CP-element group 64: 	75 
    -- CP-element group 64: 	80 
    -- CP-element group 64: 	85 
    -- CP-element group 64: 	90 
    -- CP-element group 64: 	95 
    -- CP-element group 64:  members (30) 
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/word_access_complete/$exit
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/word_access_complete/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/word_access_complete/word_0/ca
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/ptr_deref_940_Merge/$entry
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/ptr_deref_940_Merge/$exit
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/ptr_deref_940_Merge/merge_req
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_940_Update/ptr_deref_940_Merge/merge_ack
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_Sample/rr
      -- 
    ca_2684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_940_load_0_ack_1, ack => sendB_CP_2093_elements(64)); -- 
    rr_2697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(64), ack => type_cast_950_inst_req_0); -- 
    rr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(64), ack => type_cast_971_inst_req_0); -- 
    rr_2825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(64), ack => type_cast_992_inst_req_0); -- 
    rr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(64), ack => type_cast_1013_inst_req_0); -- 
    rr_2953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(64), ack => type_cast_1034_inst_req_0); -- 
    rr_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(64), ack => type_cast_1055_inst_req_0); -- 
    rr_3081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(64), ack => type_cast_1076_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_Sample/ra
      -- 
    ra_2698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_950_inst_ack_0, ack => sendB_CP_2093_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	56 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_950_Update/ca
      -- 
    ca_2703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_950_inst_ack_1, ack => sendB_CP_2093_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	56 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/ptr_deref_960_Split/$entry
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/ptr_deref_960_Split/$exit
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/ptr_deref_960_Split/split_req
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/ptr_deref_960_Split/split_ack
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/word_access_start/$entry
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/word_access_start/word_0/$entry
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/word_access_start/word_0/rr
      -- 
    rr_2741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(67), ack => ptr_deref_960_store_0_req_0); -- 
    sendB_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(56) & sendB_CP_2093_elements(66);
      gj_sendB_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	100 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/word_access_start/$exit
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/word_access_start/word_0/$exit
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Sample/word_access_start/word_0/ra
      -- 
    ra_2742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_store_0_ack_0, ack => sendB_CP_2093_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	56 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	106 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Update/word_access_complete/$exit
      -- CP-element group 69: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Update/word_access_complete/word_0/$exit
      -- CP-element group 69: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_Update/word_access_complete/word_0/ca
      -- 
    ca_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_960_store_0_ack_1, ack => sendB_CP_2093_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	64 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_Sample/ra
      -- 
    ra_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_971_inst_ack_0, ack => sendB_CP_2093_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	56 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_971_Update/ca
      -- 
    ca_2767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_971_inst_ack_1, ack => sendB_CP_2093_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	56 
    -- CP-element group 72: 	71 
    -- CP-element group 72: 	100 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (9) 
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/word_access_start/word_0/rr
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/word_access_start/word_0/$entry
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/word_access_start/$entry
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/ptr_deref_981_Split/split_ack
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/ptr_deref_981_Split/split_req
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/ptr_deref_981_Split/$exit
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/ptr_deref_981_Split/$entry
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_sample_start_
      -- 
    rr_2805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(72), ack => ptr_deref_981_store_0_req_0); -- 
    sendB_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(56) & sendB_CP_2093_elements(71) & sendB_CP_2093_elements(100);
      gj_sendB_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	101 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/word_access_start/word_0/ra
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/word_access_start/word_0/$exit
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/word_access_start/$exit
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_sample_completed_
      -- 
    ra_2806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_981_store_0_ack_0, ack => sendB_CP_2093_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	56 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	106 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Update/word_access_complete/$exit
      -- CP-element group 74: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Update/word_access_complete/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_Update/word_access_complete/word_0/ca
      -- 
    ca_2817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_981_store_0_ack_1, ack => sendB_CP_2093_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	64 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_sample_completed_
      -- 
    ra_2826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_992_inst_ack_0, ack => sendB_CP_2093_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	56 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_992_Update/ca
      -- 
    ca_2831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_992_inst_ack_1, ack => sendB_CP_2093_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	56 
    -- CP-element group 77: 	76 
    -- CP-element group 77: 	101 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/ptr_deref_1002_Split/$exit
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/ptr_deref_1002_Split/$entry
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/ptr_deref_1002_Split/split_req
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/ptr_deref_1002_Split/split_ack
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/$entry
      -- 
    rr_2869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(77), ack => ptr_deref_1002_store_0_req_0); -- 
    sendB_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(56) & sendB_CP_2093_elements(76) & sendB_CP_2093_elements(101);
      gj_sendB_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	102 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/word_access_start/$exit
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/word_access_start/word_0/$exit
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Sample/word_access_start/word_0/ra
      -- 
    ra_2870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_store_0_ack_0, ack => sendB_CP_2093_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	56 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	106 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Update/word_access_complete/word_0/ca
      -- CP-element group 79: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Update/word_access_complete/word_0/$exit
      -- CP-element group 79: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Update/word_access_complete/$exit
      -- CP-element group 79: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_Update/$exit
      -- 
    ca_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1002_store_0_ack_1, ack => sendB_CP_2093_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	64 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_Sample/ra
      -- CP-element group 80: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_sample_completed_
      -- 
    ra_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1013_inst_ack_0, ack => sendB_CP_2093_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	56 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1013_update_completed_
      -- 
    ca_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1013_inst_ack_1, ack => sendB_CP_2093_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	56 
    -- CP-element group 82: 	81 
    -- CP-element group 82: 	102 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (9) 
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/ptr_deref_1023_Split/$entry
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/word_access_start/word_0/rr
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/word_access_start/word_0/$entry
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/word_access_start/$entry
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/ptr_deref_1023_Split/split_ack
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/ptr_deref_1023_Split/split_req
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/ptr_deref_1023_Split/$exit
      -- 
    rr_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(82), ack => ptr_deref_1023_store_0_req_0); -- 
    sendB_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(56) & sendB_CP_2093_elements(81) & sendB_CP_2093_elements(102);
      gj_sendB_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	103 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/word_access_start/word_0/ra
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/word_access_start/word_0/$exit
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Sample/word_access_start/$exit
      -- 
    ra_2934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1023_store_0_ack_0, ack => sendB_CP_2093_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	56 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	106 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Update/word_access_complete/word_0/ca
      -- CP-element group 84: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Update/word_access_complete/word_0/$exit
      -- CP-element group 84: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Update/word_access_complete/$exit
      -- CP-element group 84: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_Update/$exit
      -- 
    ca_2945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1023_store_0_ack_1, ack => sendB_CP_2093_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	64 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_Sample/ra
      -- 
    ra_2954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1034_inst_ack_0, ack => sendB_CP_2093_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	56 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1034_Update/$exit
      -- 
    ca_2959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1034_inst_ack_1, ack => sendB_CP_2093_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	56 
    -- CP-element group 87: 	86 
    -- CP-element group 87: 	103 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/ptr_deref_1044_Split/$entry
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/ptr_deref_1044_Split/$exit
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/ptr_deref_1044_Split/split_req
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/ptr_deref_1044_Split/split_ack
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/word_access_start/$entry
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/word_access_start/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/word_access_start/word_0/rr
      -- 
    rr_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(87), ack => ptr_deref_1044_store_0_req_0); -- 
    sendB_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(56) & sendB_CP_2093_elements(86) & sendB_CP_2093_elements(103);
      gj_sendB_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	104 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/word_access_start/$exit
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/word_access_start/word_0/$exit
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Sample/word_access_start/word_0/ra
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_sample_completed_
      -- 
    ra_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1044_store_0_ack_0, ack => sendB_CP_2093_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	56 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	106 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Update/word_access_complete/word_0/ca
      -- CP-element group 89: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Update/word_access_complete/word_0/$exit
      -- CP-element group 89: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Update/word_access_complete/$exit
      -- CP-element group 89: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_Update/$exit
      -- 
    ca_3009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1044_store_0_ack_1, ack => sendB_CP_2093_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	64 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_sample_completed_
      -- 
    ra_3018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_0, ack => sendB_CP_2093_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	56 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1055_update_completed_
      -- 
    ca_3023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1055_inst_ack_1, ack => sendB_CP_2093_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	56 
    -- CP-element group 92: 	91 
    -- CP-element group 92: 	104 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/ptr_deref_1065_Split/$entry
      -- CP-element group 92: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/ptr_deref_1065_Split/$exit
      -- CP-element group 92: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/ptr_deref_1065_Split/split_req
      -- CP-element group 92: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/ptr_deref_1065_Split/split_ack
      -- CP-element group 92: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/word_access_start/$entry
      -- CP-element group 92: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/word_access_start/word_0/rr
      -- CP-element group 92: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/word_access_start/word_0/$entry
      -- 
    rr_3061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(92), ack => ptr_deref_1065_store_0_req_0); -- 
    sendB_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(56) & sendB_CP_2093_elements(91) & sendB_CP_2093_elements(104);
      gj_sendB_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	105 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/word_access_start/word_0/ra
      -- CP-element group 93: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/word_access_start/word_0/$exit
      -- CP-element group 93: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Sample/word_access_start/$exit
      -- 
    ra_3062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1065_store_0_ack_0, ack => sendB_CP_2093_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	56 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	106 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Update/word_access_complete/$exit
      -- CP-element group 94: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Update/word_access_complete/word_0/ca
      -- CP-element group 94: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_Update/word_access_complete/word_0/$exit
      -- 
    ca_3073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1065_store_0_ack_1, ack => sendB_CP_2093_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	64 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_sample_completed_
      -- 
    ra_3082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1076_inst_ack_0, ack => sendB_CP_2093_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	56 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/type_cast_1076_update_completed_
      -- 
    ca_3087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1076_inst_ack_1, ack => sendB_CP_2093_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	56 
    -- CP-element group 97: 	96 
    -- CP-element group 97: 	105 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (9) 
      -- CP-element group 97: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/word_access_start/word_0/rr
      -- CP-element group 97: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/word_access_start/word_0/$entry
      -- CP-element group 97: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/word_access_start/$entry
      -- CP-element group 97: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/ptr_deref_1086_Split/split_ack
      -- CP-element group 97: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/ptr_deref_1086_Split/split_req
      -- CP-element group 97: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/ptr_deref_1086_Split/$exit
      -- CP-element group 97: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/ptr_deref_1086_Split/$entry
      -- 
    rr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(97), ack => ptr_deref_1086_store_0_req_0); -- 
    sendB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(56) & sendB_CP_2093_elements(96) & sendB_CP_2093_elements(105);
      gj_sendB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (5) 
      -- CP-element group 98: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/word_access_start/word_0/ra
      -- CP-element group 98: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/word_access_start/word_0/$exit
      -- CP-element group 98: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/word_access_start/$exit
      -- CP-element group 98: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Sample/$exit
      -- 
    ra_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1086_store_0_ack_0, ack => sendB_CP_2093_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	56 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	106 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Update/word_access_complete/$exit
      -- CP-element group 99: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Update/word_access_complete/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1086_Update/word_access_complete/word_0/ca
      -- 
    ca_3137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1086_store_0_ack_1, ack => sendB_CP_2093_elements(99)); -- 
    -- CP-element group 100:  transition  delay-element  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	68 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	72 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_960_ptr_deref_981_delay
      -- 
    -- Element group sendB_CP_2093_elements(100) is a control-delay.
    cp_element_100_delay: control_delay_element  generic map(name => " 100_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(68), ack => sendB_CP_2093_elements(100), clk => clk, reset =>reset);
    -- CP-element group 101:  transition  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	73 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	77 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_981_ptr_deref_1002_delay
      -- 
    -- Element group sendB_CP_2093_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(73), ack => sendB_CP_2093_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  transition  delay-element  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	78 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	82 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1002_ptr_deref_1023_delay
      -- 
    -- Element group sendB_CP_2093_elements(102) is a control-delay.
    cp_element_102_delay: control_delay_element  generic map(name => " 102_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(78), ack => sendB_CP_2093_elements(102), clk => clk, reset =>reset);
    -- CP-element group 103:  transition  delay-element  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	83 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	87 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1023_ptr_deref_1044_delay
      -- 
    -- Element group sendB_CP_2093_elements(103) is a control-delay.
    cp_element_103_delay: control_delay_element  generic map(name => " 103_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(83), ack => sendB_CP_2093_elements(103), clk => clk, reset =>reset);
    -- CP-element group 104:  transition  delay-element  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	88 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	92 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1044_ptr_deref_1065_delay
      -- 
    -- Element group sendB_CP_2093_elements(104) is a control-delay.
    cp_element_104_delay: control_delay_element  generic map(name => " 104_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(88), ack => sendB_CP_2093_elements(104), clk => clk, reset =>reset);
    -- CP-element group 105:  transition  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	93 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	97 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/ptr_deref_1065_ptr_deref_1086_delay
      -- 
    -- Element group sendB_CP_2093_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(93), ack => sendB_CP_2093_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  branch  join  transition  place  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	58 
    -- CP-element group 106: 	59 
    -- CP-element group 106: 	69 
    -- CP-element group 106: 	74 
    -- CP-element group 106: 	79 
    -- CP-element group 106: 	84 
    -- CP-element group 106: 	89 
    -- CP-element group 106: 	94 
    -- CP-element group 106: 	99 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (10) 
      -- CP-element group 106: 	 branch_block_stmt_689/if_stmt_1095_eval_test/branch_req
      -- CP-element group 106: 	 branch_block_stmt_689/if_stmt_1095__entry__
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094__exit__
      -- CP-element group 106: 	 branch_block_stmt_689/if_stmt_1095_if_link/$entry
      -- CP-element group 106: 	 branch_block_stmt_689/if_stmt_1095_else_link/$entry
      -- CP-element group 106: 	 branch_block_stmt_689/if_stmt_1095_eval_test/$exit
      -- CP-element group 106: 	 branch_block_stmt_689/if_stmt_1095_eval_test/$entry
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_930_to_assign_stmt_1094/$exit
      -- CP-element group 106: 	 branch_block_stmt_689/R_cmp53x_xi_1096_place
      -- CP-element group 106: 	 branch_block_stmt_689/if_stmt_1095_dead_link/$entry
      -- 
    branch_req_3151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(106), ack => if_stmt_1095_branch_req_0); -- 
    sendB_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(58) & sendB_CP_2093_elements(59) & sendB_CP_2093_elements(69) & sendB_CP_2093_elements(74) & sendB_CP_2093_elements(79) & sendB_CP_2093_elements(84) & sendB_CP_2093_elements(89) & sendB_CP_2093_elements(94) & sendB_CP_2093_elements(99);
      gj_sendB_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  place  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	145 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_689/if_stmt_1095_if_link/$exit
      -- CP-element group 107: 	 branch_block_stmt_689/if_stmt_1095_if_link/if_choice_transition
      -- CP-element group 107: 	 branch_block_stmt_689/ifx_xthen_sendRemainingElementsx_xexit
      -- CP-element group 107: 	 branch_block_stmt_689/ifx_xthen_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 107: 	 branch_block_stmt_689/ifx_xthen_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_3156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1095_branch_ack_1, ack => sendB_CP_2093_elements(107)); -- 
    -- CP-element group 108:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	110 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (21) 
      -- CP-element group 108: 	 branch_block_stmt_689/ifx_xthen_bbx_xnphx_xi
      -- CP-element group 108: 	 branch_block_stmt_689/merge_stmt_1101__exit__
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145__entry__
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_update_start_
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_Sample/req
      -- CP-element group 108: 	 branch_block_stmt_689/if_stmt_1095_else_link/$exit
      -- CP-element group 108: 	 branch_block_stmt_689/if_stmt_1095_else_link/else_choice_transition
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/$entry
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_Update/cr
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_689/ifx_xthen_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 108: 	 branch_block_stmt_689/ifx_xthen_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 108: 	 branch_block_stmt_689/merge_stmt_1101_PhiReqMerge
      -- CP-element group 108: 	 branch_block_stmt_689/merge_stmt_1101_PhiAck/$entry
      -- CP-element group 108: 	 branch_block_stmt_689/merge_stmt_1101_PhiAck/$exit
      -- CP-element group 108: 	 branch_block_stmt_689/merge_stmt_1101_PhiAck/dummy
      -- 
    else_choice_transition_3160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1095_branch_ack_0, ack => sendB_CP_2093_elements(108)); -- 
    req_3187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(108), ack => WPIPE_maxpool_output_pipe_1137_inst_req_0); -- 
    cr_3178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(108), ack => type_cast_1104_inst_req_1); -- 
    rr_3173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(108), ack => type_cast_1104_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_Sample/$exit
      -- 
    ra_3174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_0, ack => sendB_CP_2093_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/type_cast_1104_Update/ca
      -- 
    ca_3179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_1, ack => sendB_CP_2093_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_Update/req
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_Sample/ack
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_update_start_
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_Sample/$exit
      -- 
    ack_3188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1137_inst_ack_0, ack => sendB_CP_2093_elements(111)); -- 
    req_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(111), ack => WPIPE_maxpool_output_pipe_1137_inst_req_1); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_Update/ack
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/WPIPE_maxpool_output_pipe_1137_update_completed_
      -- 
    ack_3193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1137_inst_ack_1, ack => sendB_CP_2093_elements(112)); -- 
    -- CP-element group 113:  branch  join  transition  place  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (10) 
      -- CP-element group 113: 	 branch_block_stmt_689/R_exitcondx_xi73_1147_place
      -- CP-element group 113: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145__exit__
      -- CP-element group 113: 	 branch_block_stmt_689/if_stmt_1146__entry__
      -- CP-element group 113: 	 branch_block_stmt_689/if_stmt_1146_if_link/$entry
      -- CP-element group 113: 	 branch_block_stmt_689/if_stmt_1146_dead_link/$entry
      -- CP-element group 113: 	 branch_block_stmt_689/if_stmt_1146_eval_test/$entry
      -- CP-element group 113: 	 branch_block_stmt_689/if_stmt_1146_eval_test/$exit
      -- CP-element group 113: 	 branch_block_stmt_689/assign_stmt_1105_to_assign_stmt_1145/$exit
      -- CP-element group 113: 	 branch_block_stmt_689/if_stmt_1146_eval_test/branch_req
      -- CP-element group 113: 	 branch_block_stmt_689/if_stmt_1146_else_link/$entry
      -- 
    branch_req_3201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(113), ack => if_stmt_1146_branch_req_0); -- 
    sendB_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(110) & sendB_CP_2093_elements(112);
      gj_sendB_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  place  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	145 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_689/bbx_xnphx_xi_sendRemainingElementsx_xexit
      -- CP-element group 114: 	 branch_block_stmt_689/if_stmt_1146_if_link/$exit
      -- CP-element group 114: 	 branch_block_stmt_689/if_stmt_1146_if_link/if_choice_transition
      -- CP-element group 114: 	 branch_block_stmt_689/bbx_xnphx_xi_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 114: 	 branch_block_stmt_689/bbx_xnphx_xi_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_3206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1146_branch_ack_1, ack => sendB_CP_2093_elements(114)); -- 
    -- CP-element group 115:  merge  transition  place  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	139 
    -- CP-element group 115:  members (18) 
      -- CP-element group 115: 	 branch_block_stmt_689/merge_stmt_1152__exit__
      -- CP-element group 115: 	 branch_block_stmt_689/assign_stmt_1158__entry__
      -- CP-element group 115: 	 branch_block_stmt_689/bbx_xnphx_xi_bbx_xnph
      -- CP-element group 115: 	 branch_block_stmt_689/bbx_xnph_forx_xbodyx_xforx_xbody_crit_edgex_xi
      -- CP-element group 115: 	 branch_block_stmt_689/assign_stmt_1158__exit__
      -- CP-element group 115: 	 branch_block_stmt_689/if_stmt_1146_else_link/else_choice_transition
      -- CP-element group 115: 	 branch_block_stmt_689/assign_stmt_1158/$entry
      -- CP-element group 115: 	 branch_block_stmt_689/assign_stmt_1158/$exit
      -- CP-element group 115: 	 branch_block_stmt_689/if_stmt_1146_else_link/$exit
      -- CP-element group 115: 	 branch_block_stmt_689/bbx_xnphx_xi_bbx_xnph_PhiReq/$entry
      -- CP-element group 115: 	 branch_block_stmt_689/bbx_xnphx_xi_bbx_xnph_PhiReq/$exit
      -- CP-element group 115: 	 branch_block_stmt_689/merge_stmt_1152_PhiReqMerge
      -- CP-element group 115: 	 branch_block_stmt_689/merge_stmt_1152_PhiAck/$entry
      -- CP-element group 115: 	 branch_block_stmt_689/merge_stmt_1152_PhiAck/$exit
      -- CP-element group 115: 	 branch_block_stmt_689/merge_stmt_1152_PhiAck/dummy
      -- CP-element group 115: 	 branch_block_stmt_689/bbx_xnph_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/$entry
      -- CP-element group 115: 	 branch_block_stmt_689/bbx_xnph_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/$entry
      -- CP-element group 115: 	 branch_block_stmt_689/bbx_xnph_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/$entry
      -- 
    else_choice_transition_3210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1146_branch_ack_0, ack => sendB_CP_2093_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	144 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	124 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_final_index_sum_regn_Sample/ack
      -- CP-element group 116: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_final_index_sum_regn_sample_complete
      -- CP-element group 116: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_final_index_sum_regn_Sample/$exit
      -- 
    ack_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1179_index_offset_ack_0, ack => sendB_CP_2093_elements(116)); -- 
    -- CP-element group 117:  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	144 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (11) 
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_request/req
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_base_plus_offset/sum_rename_ack
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_final_index_sum_regn_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_root_address_calculated
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_offset_calculated
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_base_plus_offset/sum_rename_req
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_base_plus_offset/$exit
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_base_plus_offset/$entry
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_final_index_sum_regn_Update/ack
      -- CP-element group 117: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_request/$entry
      -- 
    ack_3250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1179_index_offset_ack_1, ack => sendB_CP_2093_elements(117)); -- 
    req_3259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(117), ack => array_obj_ref_1179_final_reg_req_0); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_request/$exit
      -- CP-element group 118: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_request/ack
      -- 
    ack_3260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1179_final_reg_ack_0, ack => sendB_CP_2093_elements(118)); -- 
    -- CP-element group 119:  join  fork  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	144 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (24) 
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_complete/ack
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_complete/$exit
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_base_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_word_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_base_address_resized
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_base_addr_resize/$entry
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_base_addr_resize/$exit
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_base_addr_resize/base_resize_req
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_base_addr_resize/base_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_word_addrgen/$entry
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_word_addrgen/$exit
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_word_addrgen/root_register_req
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_word_addrgen/root_register_ack
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Sample/word_access_start/$entry
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Sample/word_access_start/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Sample/word_access_start/word_0/rr
      -- 
    ack_3265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1179_final_reg_ack_1, ack => sendB_CP_2093_elements(119)); -- 
    rr_3298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(119), ack => ptr_deref_1183_load_0_req_0); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Sample/word_access_start/$exit
      -- CP-element group 120: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Sample/word_access_start/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Sample/word_access_start/word_0/ra
      -- 
    ra_3299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1183_load_0_ack_0, ack => sendB_CP_2093_elements(120)); -- 
    -- CP-element group 121:  transition  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	144 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (12) 
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/word_access_complete/$exit
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/word_access_complete/word_0/$exit
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/word_access_complete/word_0/ca
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/ptr_deref_1183_Merge/$entry
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/ptr_deref_1183_Merge/$exit
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/ptr_deref_1183_Merge/merge_req
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/ptr_deref_1183_Merge/merge_ack
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_Sample/req
      -- 
    ca_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1183_load_0_ack_1, ack => sendB_CP_2093_elements(121)); -- 
    req_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(121), ack => WPIPE_maxpool_output_pipe_1185_inst_req_0); -- 
    -- CP-element group 122:  transition  input  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (6) 
      -- CP-element group 122: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_update_start_
      -- CP-element group 122: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_Sample/ack
      -- CP-element group 122: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_Update/req
      -- 
    ack_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1185_inst_ack_0, ack => sendB_CP_2093_elements(122)); -- 
    req_3328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(122), ack => WPIPE_maxpool_output_pipe_1185_inst_req_1); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/WPIPE_maxpool_output_pipe_1185_Update/ack
      -- 
    ack_3329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1185_inst_ack_1, ack => sendB_CP_2093_elements(123)); -- 
    -- CP-element group 124:  branch  join  transition  place  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	116 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (10) 
      -- CP-element group 124: 	 branch_block_stmt_689/if_stmt_1193__entry__
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192__exit__
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/$exit
      -- CP-element group 124: 	 branch_block_stmt_689/if_stmt_1193_dead_link/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/if_stmt_1193_eval_test/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/if_stmt_1193_eval_test/$exit
      -- CP-element group 124: 	 branch_block_stmt_689/if_stmt_1193_eval_test/branch_req
      -- CP-element group 124: 	 branch_block_stmt_689/R_exitcond3_1194_place
      -- CP-element group 124: 	 branch_block_stmt_689/if_stmt_1193_if_link/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/if_stmt_1193_else_link/$entry
      -- 
    branch_req_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => if_stmt_1193_branch_req_0); -- 
    sendB_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(116) & sendB_CP_2093_elements(123);
      gj_sendB_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  place  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	145 
    -- CP-element group 125:  members (13) 
      -- CP-element group 125: 	 branch_block_stmt_689/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit
      -- CP-element group 125: 	 branch_block_stmt_689/merge_stmt_1207__exit__
      -- CP-element group 125: 	 branch_block_stmt_689/if_stmt_1193_if_link/$exit
      -- CP-element group 125: 	 branch_block_stmt_689/if_stmt_1193_if_link/if_choice_transition
      -- CP-element group 125: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xi_sendRemainingElementsx_xexitx_xloopexit
      -- CP-element group 125: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xi_sendRemainingElementsx_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xi_sendRemainingElementsx_xexitx_xloopexit_PhiReq/$exit
      -- CP-element group 125: 	 branch_block_stmt_689/merge_stmt_1207_PhiReqMerge
      -- CP-element group 125: 	 branch_block_stmt_689/merge_stmt_1207_PhiAck/$entry
      -- CP-element group 125: 	 branch_block_stmt_689/merge_stmt_1207_PhiAck/$exit
      -- CP-element group 125: 	 branch_block_stmt_689/merge_stmt_1207_PhiAck/dummy
      -- CP-element group 125: 	 branch_block_stmt_689/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_689/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_3342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1193_branch_ack_1, ack => sendB_CP_2093_elements(125)); -- 
    -- CP-element group 126:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	140 
    -- CP-element group 126: 	141 
    -- CP-element group 126:  members (24) 
      -- CP-element group 126: 	 branch_block_stmt_689/merge_stmt_1199__exit__
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi
      -- CP-element group 126: 	 branch_block_stmt_689/assign_stmt_1205__exit__
      -- CP-element group 126: 	 branch_block_stmt_689/assign_stmt_1205__entry__
      -- CP-element group 126: 	 branch_block_stmt_689/if_stmt_1193_else_link/$exit
      -- CP-element group 126: 	 branch_block_stmt_689/if_stmt_1193_else_link/else_choice_transition
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xi_forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge
      -- CP-element group 126: 	 branch_block_stmt_689/assign_stmt_1205/$entry
      -- CP-element group 126: 	 branch_block_stmt_689/assign_stmt_1205/$exit
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/$entry
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/$entry
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/$entry
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/$entry
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/$entry
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Sample/rr
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Update/cr
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xi_forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_PhiReq/$entry
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xi_forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_PhiReq/$exit
      -- CP-element group 126: 	 branch_block_stmt_689/merge_stmt_1199_PhiReqMerge
      -- CP-element group 126: 	 branch_block_stmt_689/merge_stmt_1199_PhiAck/$entry
      -- CP-element group 126: 	 branch_block_stmt_689/merge_stmt_1199_PhiAck/$exit
      -- CP-element group 126: 	 branch_block_stmt_689/merge_stmt_1199_PhiAck/dummy
      -- 
    else_choice_transition_3346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1193_branch_ack_0, ack => sendB_CP_2093_elements(126)); -- 
    rr_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(126), ack => type_cast_1164_inst_req_0); -- 
    cr_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(126), ack => type_cast_1164_inst_req_1); -- 
    -- CP-element group 127:  transition  output  delay-element  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	4 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	131 
    -- CP-element group 127:  members (5) 
      -- CP-element group 127: 	 branch_block_stmt_689/bbx_xnph78_forx_xbody_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_689/bbx_xnph78_forx_xbody_PhiReq/phi_stmt_752/$exit
      -- CP-element group 127: 	 branch_block_stmt_689/bbx_xnph78_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/$exit
      -- CP-element group 127: 	 branch_block_stmt_689/bbx_xnph78_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_756_konst_delay_trans
      -- CP-element group 127: 	 branch_block_stmt_689/bbx_xnph78_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_req
      -- 
    phi_stmt_752_req_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_752_req_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(127), ack => phi_stmt_752_req_0); -- 
    -- Element group sendB_CP_2093_elements(127) is a control-delay.
    cp_element_127_delay: control_delay_element  generic map(name => " 127_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(4), ack => sendB_CP_2093_elements(127), clk => clk, reset =>reset);
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	52 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/SplitProtocol/Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/SplitProtocol/Sample/ra
      -- 
    ra_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_758_inst_ack_0, ack => sendB_CP_2093_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	52 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/SplitProtocol/Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/SplitProtocol/Update/ca
      -- 
    ca_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_758_inst_ack_1, ack => sendB_CP_2093_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (6) 
      -- CP-element group 130: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/$exit
      -- CP-element group 130: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/$exit
      -- CP-element group 130: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/$exit
      -- CP-element group 130: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_sources/type_cast_758/SplitProtocol/$exit
      -- CP-element group 130: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_752/phi_stmt_752_req
      -- 
    phi_stmt_752_req_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_752_req_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(130), ack => phi_stmt_752_req_1); -- 
    sendB_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(128) & sendB_CP_2093_elements(129);
      gj_sendB_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  merge  transition  place  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	127 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_689/merge_stmt_751_PhiReqMerge
      -- CP-element group 131: 	 branch_block_stmt_689/merge_stmt_751_PhiAck/$entry
      -- 
    sendB_CP_2093_elements(131) <= OrReduce(sendB_CP_2093_elements(127) & sendB_CP_2093_elements(130));
    -- CP-element group 132:  fork  transition  place  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	5 
    -- CP-element group 132: 	6 
    -- CP-element group 132: 	8 
    -- CP-element group 132: 	10 
    -- CP-element group 132: 	12 
    -- CP-element group 132: 	14 
    -- CP-element group 132: 	16 
    -- CP-element group 132: 	18 
    -- CP-element group 132: 	20 
    -- CP-element group 132: 	22 
    -- CP-element group 132: 	24 
    -- CP-element group 132: 	26 
    -- CP-element group 132:  members (53) 
      -- CP-element group 132: 	 branch_block_stmt_689/merge_stmt_751__exit__
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879__entry__
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_update_start_
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_resized_1
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_scaled_1
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_computed_1
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_resize_1/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_resize_1/$exit
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_resize_1/index_resize_req
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_resize_1/index_resize_ack
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_scale_1/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_scale_1/$exit
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_scale_1/scale_rename_req
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_index_scale_1/scale_rename_ack
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_final_index_sum_regn_update_start
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_final_index_sum_regn_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_final_index_sum_regn_Sample/req
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_final_index_sum_regn_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/array_obj_ref_764_final_index_sum_regn_Update/req
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_complete/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/addr_of_765_complete/req
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_update_start_
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/word_access_complete/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/word_access_complete/word_0/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/ptr_deref_769_Update/word_access_complete/word_0/cr
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_update_start_
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_773_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_update_start_
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_783_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_update_start_
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_793_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_update_start_
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_803_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_update_start_
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_813_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_update_start_
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_823_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_update_start_
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_833_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_update_start_
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_689/assign_stmt_766_to_assign_stmt_879/type_cast_843_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_689/merge_stmt_751_PhiAck/$exit
      -- CP-element group 132: 	 branch_block_stmt_689/merge_stmt_751_PhiAck/phi_stmt_752_ack
      -- 
    phi_stmt_752_ack_3405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_752_ack_0, ack => sendB_CP_2093_elements(132)); -- 
    req_2223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => array_obj_ref_764_index_offset_req_0); -- 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => array_obj_ref_764_index_offset_req_1); -- 
    req_2243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => addr_of_765_final_reg_req_1); -- 
    cr_2288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => ptr_deref_769_load_0_req_1); -- 
    cr_2307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => type_cast_773_inst_req_1); -- 
    cr_2321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => type_cast_783_inst_req_1); -- 
    cr_2335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => type_cast_793_inst_req_1); -- 
    cr_2349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => type_cast_803_inst_req_1); -- 
    cr_2363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => type_cast_813_inst_req_1); -- 
    cr_2377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => type_cast_823_inst_req_1); -- 
    cr_2391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => type_cast_833_inst_req_1); -- 
    cr_2405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(132), ack => type_cast_843_inst_req_1); -- 
    -- CP-element group 133:  transition  output  delay-element  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	2 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	137 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/$exit
      -- CP-element group 133: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_900/$exit
      -- CP-element group 133: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/$exit
      -- CP-element group 133: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_906_konst_delay_trans
      -- CP-element group 133: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_req
      -- 
    phi_stmt_900_req_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_900_req_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(133), ack => phi_stmt_900_req_1); -- 
    -- Element group sendB_CP_2093_elements(133) is a control-delay.
    cp_element_133_delay: control_delay_element  generic map(name => " 133_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(2), ack => sendB_CP_2093_elements(133), clk => clk, reset =>reset);
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	54 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/SplitProtocol/Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/SplitProtocol/Sample/ra
      -- 
    ra_3448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_0, ack => sendB_CP_2093_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	54 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/SplitProtocol/Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/SplitProtocol/Update/ca
      -- 
    ca_3453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_903_inst_ack_1, ack => sendB_CP_2093_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (6) 
      -- CP-element group 136: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 136: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/$exit
      -- CP-element group 136: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/$exit
      -- CP-element group 136: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/$exit
      -- CP-element group 136: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_sources/type_cast_903/SplitProtocol/$exit
      -- CP-element group 136: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_900/phi_stmt_900_req
      -- 
    phi_stmt_900_req_3454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_900_req_3454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(136), ack => phi_stmt_900_req_0); -- 
    sendB_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(134) & sendB_CP_2093_elements(135);
      gj_sendB_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  merge  transition  place  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	133 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (2) 
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_899_PhiReqMerge
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_899_PhiAck/$entry
      -- 
    sendB_CP_2093_elements(137) <= OrReduce(sendB_CP_2093_elements(133) & sendB_CP_2093_elements(136));
    -- CP-element group 138:  branch  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	55 
    -- CP-element group 138: 	56 
    -- CP-element group 138:  members (15) 
      -- CP-element group 138: 	 branch_block_stmt_689/assign_stmt_913_to_assign_stmt_919__exit__
      -- CP-element group 138: 	 branch_block_stmt_689/assign_stmt_913_to_assign_stmt_919__entry__
      -- CP-element group 138: 	 branch_block_stmt_689/if_stmt_920__entry__
      -- CP-element group 138: 	 branch_block_stmt_689/merge_stmt_899__exit__
      -- CP-element group 138: 	 branch_block_stmt_689/assign_stmt_913_to_assign_stmt_919/$entry
      -- CP-element group 138: 	 branch_block_stmt_689/assign_stmt_913_to_assign_stmt_919/$exit
      -- CP-element group 138: 	 branch_block_stmt_689/if_stmt_920_dead_link/$entry
      -- CP-element group 138: 	 branch_block_stmt_689/if_stmt_920_eval_test/$entry
      -- CP-element group 138: 	 branch_block_stmt_689/if_stmt_920_eval_test/$exit
      -- CP-element group 138: 	 branch_block_stmt_689/if_stmt_920_eval_test/branch_req
      -- CP-element group 138: 	 branch_block_stmt_689/R_tobool_921_place
      -- CP-element group 138: 	 branch_block_stmt_689/if_stmt_920_if_link/$entry
      -- CP-element group 138: 	 branch_block_stmt_689/if_stmt_920_else_link/$entry
      -- CP-element group 138: 	 branch_block_stmt_689/merge_stmt_899_PhiAck/$exit
      -- CP-element group 138: 	 branch_block_stmt_689/merge_stmt_899_PhiAck/phi_stmt_900_ack
      -- 
    phi_stmt_900_ack_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_900_ack_0, ack => sendB_CP_2093_elements(138)); -- 
    branch_req_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(138), ack => if_stmt_920_branch_req_0); -- 
    -- CP-element group 139:  transition  output  delay-element  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	115 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	143 
    -- CP-element group 139:  members (5) 
      -- CP-element group 139: 	 branch_block_stmt_689/bbx_xnph_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/$exit
      -- CP-element group 139: 	 branch_block_stmt_689/bbx_xnph_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/$exit
      -- CP-element group 139: 	 branch_block_stmt_689/bbx_xnph_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/$exit
      -- CP-element group 139: 	 branch_block_stmt_689/bbx_xnph_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1167_konst_delay_trans
      -- CP-element group 139: 	 branch_block_stmt_689/bbx_xnph_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_req
      -- 
    phi_stmt_1161_req_3506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1161_req_3506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(139), ack => phi_stmt_1161_req_1); -- 
    -- Element group sendB_CP_2093_elements(139) is a control-delay.
    cp_element_139_delay: control_delay_element  generic map(name => " 139_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(115), ack => sendB_CP_2093_elements(139), clk => clk, reset =>reset);
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	126 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Sample/ra
      -- 
    ra_3526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1164_inst_ack_0, ack => sendB_CP_2093_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	126 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/Update/ca
      -- 
    ca_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1164_inst_ack_1, ack => sendB_CP_2093_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (6) 
      -- CP-element group 142: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/$exit
      -- CP-element group 142: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/$exit
      -- CP-element group 142: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/$exit
      -- CP-element group 142: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/$exit
      -- CP-element group 142: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_sources/type_cast_1164/SplitProtocol/$exit
      -- CP-element group 142: 	 branch_block_stmt_689/forx_xbodyx_xforx_xbody_crit_edgex_xix_xforx_xbodyx_xforx_xbody_crit_edgex_xi_crit_edge_forx_xbodyx_xforx_xbody_crit_edgex_xi_PhiReq/phi_stmt_1161/phi_stmt_1161_req
      -- 
    phi_stmt_1161_req_3532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1161_req_3532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(142), ack => phi_stmt_1161_req_0); -- 
    sendB_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(140) & sendB_CP_2093_elements(141);
      gj_sendB_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  merge  transition  place  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	139 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (2) 
      -- CP-element group 143: 	 branch_block_stmt_689/merge_stmt_1160_PhiReqMerge
      -- CP-element group 143: 	 branch_block_stmt_689/merge_stmt_1160_PhiAck/$entry
      -- 
    sendB_CP_2093_elements(143) <= OrReduce(sendB_CP_2093_elements(139) & sendB_CP_2093_elements(142));
    -- CP-element group 144:  fork  transition  place  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	116 
    -- CP-element group 144: 	117 
    -- CP-element group 144: 	119 
    -- CP-element group 144: 	121 
    -- CP-element group 144:  members (29) 
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192__entry__
      -- CP-element group 144: 	 branch_block_stmt_689/merge_stmt_1160__exit__
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_complete/req
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_complete/$entry
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_resized_1
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_scaled_1
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_computed_1
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_resize_1/$entry
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_resize_1/$exit
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_resize_1/index_resize_req
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_resize_1/index_resize_ack
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_update_start_
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_final_index_sum_regn_update_start
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_final_index_sum_regn_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_final_index_sum_regn_Sample/req
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_scale_1/$entry
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_scale_1/$exit
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_scale_1/scale_rename_req
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_final_index_sum_regn_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_index_scale_1/scale_rename_ack
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/$entry
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/array_obj_ref_1179_final_index_sum_regn_Update/req
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_update_start_
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/word_access_complete/$entry
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/word_access_complete/word_0/$entry
      -- CP-element group 144: 	 branch_block_stmt_689/assign_stmt_1174_to_assign_stmt_1192/ptr_deref_1183_Update/word_access_complete/word_0/cr
      -- CP-element group 144: 	 branch_block_stmt_689/merge_stmt_1160_PhiAck/$exit
      -- CP-element group 144: 	 branch_block_stmt_689/merge_stmt_1160_PhiAck/phi_stmt_1161_ack
      -- 
    phi_stmt_1161_ack_3537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1161_ack_0, ack => sendB_CP_2093_elements(144)); -- 
    req_3264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(144), ack => array_obj_ref_1179_final_reg_req_1); -- 
    req_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(144), ack => array_obj_ref_1179_index_offset_req_0); -- 
    req_3249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(144), ack => array_obj_ref_1179_index_offset_req_1); -- 
    cr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(144), ack => ptr_deref_1183_load_0_req_1); -- 
    -- CP-element group 145:  merge  transition  place  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	55 
    -- CP-element group 145: 	107 
    -- CP-element group 145: 	114 
    -- CP-element group 145: 	125 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (16) 
      -- CP-element group 145: 	 branch_block_stmt_689/merge_stmt_1211__exit__
      -- CP-element group 145: 	 branch_block_stmt_689/merge_stmt_1209__exit__
      -- CP-element group 145: 	 branch_block_stmt_689/return__
      -- CP-element group 145: 	 $exit
      -- CP-element group 145: 	 branch_block_stmt_689/$exit
      -- CP-element group 145: 	 branch_block_stmt_689/branch_block_stmt_689__exit__
      -- CP-element group 145: 	 branch_block_stmt_689/merge_stmt_1209_PhiReqMerge
      -- CP-element group 145: 	 branch_block_stmt_689/merge_stmt_1209_PhiAck/$entry
      -- CP-element group 145: 	 branch_block_stmt_689/merge_stmt_1209_PhiAck/$exit
      -- CP-element group 145: 	 branch_block_stmt_689/merge_stmt_1209_PhiAck/dummy
      -- CP-element group 145: 	 branch_block_stmt_689/return___PhiReq/$entry
      -- CP-element group 145: 	 branch_block_stmt_689/return___PhiReq/$exit
      -- CP-element group 145: 	 branch_block_stmt_689/merge_stmt_1211_PhiReqMerge
      -- CP-element group 145: 	 branch_block_stmt_689/merge_stmt_1211_PhiAck/$entry
      -- CP-element group 145: 	 branch_block_stmt_689/merge_stmt_1211_PhiAck/$exit
      -- CP-element group 145: 	 branch_block_stmt_689/merge_stmt_1211_PhiAck/dummy
      -- 
    sendB_CP_2093_elements(145) <= OrReduce(sendB_CP_2093_elements(55) & sendB_CP_2093_elements(107) & sendB_CP_2093_elements(114) & sendB_CP_2093_elements(125));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar81_763_resized : std_logic_vector(13 downto 0);
    signal R_indvar81_763_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_934_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_934_scaled : std_logic_vector(13 downto 0);
    signal R_tmp_1178_resized : std_logic_vector(2 downto 0);
    signal R_tmp_1178_scaled : std_logic_vector(2 downto 0);
    signal and68_913 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1179_constant_part_of_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1179_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1179_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1179_offset_scale_factor_1 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1179_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1179_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_764_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_764_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_764_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_764_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_764_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_764_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_935_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_935_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_935_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_935_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_935_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_935_root_address : std_logic_vector(13 downto 0);
    signal arrayidx11x_xi_979 : std_logic_vector(31 downto 0);
    signal arrayidx17x_xi_1000 : std_logic_vector(31 downto 0);
    signal arrayidx23x_xi_1021 : std_logic_vector(31 downto 0);
    signal arrayidx29x_xi_1042 : std_logic_vector(31 downto 0);
    signal arrayidx35x_xi_1063 : std_logic_vector(31 downto 0);
    signal arrayidx41x_xi_1084 : std_logic_vector(31 downto 0);
    signal arrayidx49x_xphix_xtransx_xinsertx_xi_1180 : std_logic_vector(31 downto 0);
    signal arrayidx5x_xi_958 : std_logic_vector(31 downto 0);
    signal arrayidx_766 : std_logic_vector(31 downto 0);
    signal arrayidxx_xi_937 : std_logic_vector(31 downto 0);
    signal cmp53x_xi_1094 : std_logic_vector(0 downto 0);
    signal cmp76_701 : std_logic_vector(0 downto 0);
    signal conv10x_xi_972 : std_logic_vector(7 downto 0);
    signal conv12_784 : std_logic_vector(7 downto 0);
    signal conv16x_xi_993 : std_logic_vector(7 downto 0);
    signal conv18_794 : std_logic_vector(7 downto 0);
    signal conv22x_xi_1014 : std_logic_vector(7 downto 0);
    signal conv24_804 : std_logic_vector(7 downto 0);
    signal conv28x_xi_1035 : std_logic_vector(7 downto 0);
    signal conv30_814 : std_logic_vector(7 downto 0);
    signal conv34x_xi_1056 : std_logic_vector(7 downto 0);
    signal conv36_824 : std_logic_vector(7 downto 0);
    signal conv40x_xi_1077 : std_logic_vector(7 downto 0);
    signal conv42_834 : std_logic_vector(7 downto 0);
    signal conv48_844 : std_logic_vector(7 downto 0);
    signal conv72_930 : std_logic_vector(7 downto 0);
    signal conv_774 : std_logic_vector(7 downto 0);
    signal convx_xi_951 : std_logic_vector(7 downto 0);
    signal exitcond3_1192 : std_logic_vector(0 downto 0);
    signal exitcond_879 : std_logic_vector(0 downto 0);
    signal exitcondx_xi73_1145 : std_logic_vector(0 downto 0);
    signal iNsTr_30_1123 : std_logic_vector(63 downto 0);
    signal indvar1_1161 : std_logic_vector(63 downto 0);
    signal indvar81_752 : std_logic_vector(63 downto 0);
    signal indvarx_xnext82_874 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1205 : std_logic_vector(63 downto 0);
    signal ix_x0x_xlcssa_900 : std_logic_vector(63 downto 0);
    signal out_datax_xi_695 : std_logic_vector(31 downto 0);
    signal phitmp_897 : std_logic_vector(63 downto 0);
    signal ptr_deref_1002_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1002_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1002_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1002_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1002_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1002_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1023_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1023_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1023_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1023_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1023_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1023_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1044_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1044_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1044_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1044_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1044_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1044_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1065_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1065_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1065_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1065_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1065_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1065_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1086_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1086_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1086_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1086_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1086_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1086_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1183_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1183_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1183_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1183_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1183_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_769_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_769_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_769_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_769_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_769_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_940_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_940_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_940_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_940_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_940_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_960_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_960_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_960_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_960_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_960_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_960_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_981_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_981_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_981_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_981_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_981_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_981_word_offset_0 : std_logic_vector(2 downto 0);
    signal shr13x_xi_989 : std_logic_vector(63 downto 0);
    signal shr15_790 : std_logic_vector(63 downto 0);
    signal shr19x_xi_1010 : std_logic_vector(63 downto 0);
    signal shr21_800 : std_logic_vector(63 downto 0);
    signal shr25x_xi_1031 : std_logic_vector(63 downto 0);
    signal shr27_810 : std_logic_vector(63 downto 0);
    signal shr31x_xi_1052 : std_logic_vector(63 downto 0);
    signal shr33_820 : std_logic_vector(63 downto 0);
    signal shr37x_xi_1073 : std_logic_vector(63 downto 0);
    signal shr39_830 : std_logic_vector(63 downto 0);
    signal shr45_840 : std_logic_vector(63 downto 0);
    signal shr7x_xi_968 : std_logic_vector(63 downto 0);
    signal shr9_780 : std_logic_vector(63 downto 0);
    signal shr_714 : std_logic_vector(31 downto 0);
    signal shrx_xi_947 : std_logic_vector(63 downto 0);
    signal tmp1x_xi_941 : std_logic_vector(63 downto 0);
    signal tmp2_1158 : std_logic_vector(63 downto 0);
    signal tmp4_770 : std_logic_vector(63 downto 0);
    signal tmp50x_xprex_xi_1184 : std_logic_vector(7 downto 0);
    signal tmp55x_xi_1111 : std_logic_vector(0 downto 0);
    signal tmp58x_xi_1136 : std_logic_vector(63 downto 0);
    signal tmp5_726 : std_logic_vector(0 downto 0);
    signal tmp7_739 : std_logic_vector(31 downto 0);
    signal tmp80_720 : std_logic_vector(0 downto 0);
    signal tmp8_743 : std_logic_vector(63 downto 0);
    signal tmp9_749 : std_logic_vector(63 downto 0);
    signal tmp_1174 : std_logic_vector(63 downto 0);
    signal tmpx_xi_1105 : std_logic_vector(63 downto 0);
    signal tmpx_xopx_xi_1117 : std_logic_vector(63 downto 0);
    signal tobool_919 : std_logic_vector(0 downto 0);
    signal type_cast_1008_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1029_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1050_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1071_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1092_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1109_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1115_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1121_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1127_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1134_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1143_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1156_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1164_wire : std_logic_vector(63 downto 0);
    signal type_cast_1167_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1172_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1203_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_699_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_712_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_718_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_724_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_731_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_737_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_747_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_758_wire : std_logic_vector(63 downto 0);
    signal type_cast_778_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_788_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_798_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_808_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_818_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_828_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_838_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_872_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_903_wire : std_logic_vector(63 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_911_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_917_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_945_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_966_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_987_wire_constant : std_logic_vector(63 downto 0);
    signal umax6_733 : std_logic_vector(31 downto 0);
    signal umax_893 : std_logic_vector(31 downto 0);
    signal xx_xopx_xi_1129 : std_logic_vector(63 downto 0);
    signal xxsendBxxbodyxxout_datax_xi_alloc_base_address : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    array_obj_ref_1179_constant_part_of_offset <= "000";
    array_obj_ref_1179_offset_scale_factor_0 <= "111";
    array_obj_ref_1179_offset_scale_factor_1 <= "001";
    array_obj_ref_1179_resized_base_address <= "000";
    array_obj_ref_764_constant_part_of_offset <= "00000000000000";
    array_obj_ref_764_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_764_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_764_resized_base_address <= "00000000000000";
    array_obj_ref_935_constant_part_of_offset <= "00000000000000";
    array_obj_ref_935_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_935_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_935_resized_base_address <= "00000000000000";
    arrayidx11x_xi_979 <= "00000000000000000000000000000101";
    arrayidx17x_xi_1000 <= "00000000000000000000000000000100";
    arrayidx23x_xi_1021 <= "00000000000000000000000000000011";
    arrayidx29x_xi_1042 <= "00000000000000000000000000000010";
    arrayidx35x_xi_1063 <= "00000000000000000000000000000001";
    arrayidx41x_xi_1084 <= "00000000000000000000000000000000";
    arrayidx5x_xi_958 <= "00000000000000000000000000000110";
    out_datax_xi_695 <= "00000000000000000000000000000000";
    ptr_deref_1002_word_offset_0 <= "000";
    ptr_deref_1023_word_offset_0 <= "000";
    ptr_deref_1044_word_offset_0 <= "000";
    ptr_deref_1065_word_offset_0 <= "000";
    ptr_deref_1086_word_offset_0 <= "000";
    ptr_deref_1183_word_offset_0 <= "000";
    ptr_deref_769_word_offset_0 <= "00000000000000";
    ptr_deref_940_word_offset_0 <= "00000000000000";
    ptr_deref_960_word_offset_0 <= "000";
    ptr_deref_981_word_offset_0 <= "000";
    type_cast_1008_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1029_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1050_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1071_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1092_wire_constant <= "00000000";
    type_cast_1109_wire_constant <= "00000001";
    type_cast_1115_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_1121_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_1127_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1134_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1143_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1156_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111110";
    type_cast_1167_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1172_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1203_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_699_wire_constant <= "00000000000000000000000000000111";
    type_cast_712_wire_constant <= "00000000000000000000000000000011";
    type_cast_718_wire_constant <= "00000000000000000000000000000001";
    type_cast_724_wire_constant <= "00000000000000000000000000000001";
    type_cast_731_wire_constant <= "00000000000000000000000000000001";
    type_cast_737_wire_constant <= "11111111111111111111111111111111";
    type_cast_747_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_756_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_778_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_788_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_798_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_808_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_818_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_828_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_838_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_872_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_891_wire_constant <= "00000000000000000000000000000001";
    type_cast_906_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_911_wire_constant <= "00000000000000000000000000000111";
    type_cast_917_wire_constant <= "00000000000000000000000000000000";
    type_cast_945_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_966_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_987_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    xxsendBxxbodyxxout_datax_xi_alloc_base_address <= "000";
    phi_stmt_1161: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1164_wire & type_cast_1167_wire_constant;
      req <= phi_stmt_1161_req_0 & phi_stmt_1161_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1161",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1161_ack_0,
          idata => idata,
          odata => indvar1_1161,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1161
    phi_stmt_752: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_756_wire_constant & type_cast_758_wire;
      req <= phi_stmt_752_req_0 & phi_stmt_752_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_752",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_752_ack_0,
          idata => idata,
          odata => indvar81_752,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_752
    phi_stmt_900: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_903_wire & type_cast_906_wire_constant;
      req <= phi_stmt_900_req_0 & phi_stmt_900_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_900",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_900_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_900,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_900
    -- flow-through select operator MUX_1135_inst
    tmp58x_xi_1136 <= xx_xopx_xi_1129 when (tmp55x_xi_1111(0) /=  '0') else type_cast_1134_wire_constant;
    -- flow-through select operator MUX_732_inst
    umax6_733 <= shr_714 when (tmp5_726(0) /=  '0') else type_cast_731_wire_constant;
    -- flow-through select operator MUX_892_inst
    umax_893 <= shr_714 when (tmp80_720(0) /=  '0') else type_cast_891_wire_constant;
    addr_of_765_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_765_final_reg_req_0;
      addr_of_765_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_765_final_reg_req_1;
      addr_of_765_final_reg_ack_1<= rack(0);
      addr_of_765_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_765_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_764_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_766,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_936_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_936_final_reg_req_0;
      addr_of_936_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_936_final_reg_req_1;
      addr_of_936_final_reg_ack_1<= rack(0);
      addr_of_936_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_936_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_935_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidxx_xi_937,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    array_obj_ref_1179_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= array_obj_ref_1179_final_reg_req_0;
      array_obj_ref_1179_final_reg_ack_0<= wack(0);
      rreq(0) <= array_obj_ref_1179_final_reg_req_1;
      array_obj_ref_1179_final_reg_ack_1<= rack(0);
      array_obj_ref_1179_final_reg : InterlockBuffer generic map ( -- 
        name => "array_obj_ref_1179_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1179_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx49x_xphix_xtransx_xinsertx_xi_1180,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1013_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1013_inst_req_0;
      type_cast_1013_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1013_inst_req_1;
      type_cast_1013_inst_ack_1<= rack(0);
      type_cast_1013_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1013_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr19x_xi_1010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22x_xi_1014,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1034_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1034_inst_req_0;
      type_cast_1034_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1034_inst_req_1;
      type_cast_1034_inst_ack_1<= rack(0);
      type_cast_1034_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1034_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr25x_xi_1031,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28x_xi_1035,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1055_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1055_inst_req_0;
      type_cast_1055_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1055_inst_req_1;
      type_cast_1055_inst_ack_1<= rack(0);
      type_cast_1055_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1055_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr31x_xi_1052,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34x_xi_1056,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1076_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1076_inst_req_0;
      type_cast_1076_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1076_inst_req_1;
      type_cast_1076_inst_ack_1<= rack(0);
      type_cast_1076_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1076_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr37x_xi_1073,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv40x_xi_1077,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1104_inst_req_0;
      type_cast_1104_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1104_inst_req_1;
      type_cast_1104_inst_ack_1<= rack(0);
      type_cast_1104_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1104_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => and68_913,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmpx_xi_1105,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1164_inst_req_0;
      type_cast_1164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1164_inst_req_1;
      type_cast_1164_inst_ack_1<= rack(0);
      type_cast_1164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1205,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1164_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_742_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_742_inst_req_0;
      type_cast_742_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_742_inst_req_1;
      type_cast_742_inst_ack_1<= rack(0);
      type_cast_742_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_742_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp7_739,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp8_743,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_758_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_758_inst_req_0;
      type_cast_758_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_758_inst_req_1;
      type_cast_758_inst_ack_1<= rack(0);
      type_cast_758_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_758_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext82_874,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_758_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_773_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_773_inst_req_0;
      type_cast_773_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_773_inst_req_1;
      type_cast_773_inst_ack_1<= rack(0);
      type_cast_773_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_773_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_770,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_774,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_783_inst_req_0;
      type_cast_783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_783_inst_req_1;
      type_cast_783_inst_ack_1<= rack(0);
      type_cast_783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_783_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_793_inst_req_0;
      type_cast_793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_793_inst_req_1;
      type_cast_793_inst_ack_1<= rack(0);
      type_cast_793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_803_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_803_inst_req_0;
      type_cast_803_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_803_inst_req_1;
      type_cast_803_inst_ack_1<= rack(0);
      type_cast_803_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_803_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_800,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_804,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_813_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_813_inst_req_0;
      type_cast_813_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_813_inst_req_1;
      type_cast_813_inst_ack_1<= rack(0);
      type_cast_813_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_813_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_814,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_823_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_823_inst_req_0;
      type_cast_823_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_823_inst_req_1;
      type_cast_823_inst_ack_1<= rack(0);
      type_cast_823_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_823_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_820,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_824,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_833_inst_req_0;
      type_cast_833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_833_inst_req_1;
      type_cast_833_inst_ack_1<= rack(0);
      type_cast_833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_830,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_834,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_843_inst_req_0;
      type_cast_843_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_843_inst_req_1;
      type_cast_843_inst_ack_1<= rack(0);
      type_cast_843_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_840,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_844,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_896_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_896_inst_req_0;
      type_cast_896_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_896_inst_req_1;
      type_cast_896_inst_ack_1<= rack(0);
      type_cast_896_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_896_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => umax_893,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => phitmp_897,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_903_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_903_inst_req_0;
      type_cast_903_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_903_inst_req_1;
      type_cast_903_inst_ack_1<= rack(0);
      type_cast_903_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_903_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_897,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_903_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_929_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_929_inst_req_0;
      type_cast_929_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_929_inst_req_1;
      type_cast_929_inst_ack_1<= rack(0);
      type_cast_929_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_929_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => and68_913,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_930,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_950_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_950_inst_req_0;
      type_cast_950_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_950_inst_req_1;
      type_cast_950_inst_ack_1<= rack(0);
      type_cast_950_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_950_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shrx_xi_947,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_951,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_971_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_971_inst_req_0;
      type_cast_971_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_971_inst_req_1;
      type_cast_971_inst_ack_1<= rack(0);
      type_cast_971_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_971_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr7x_xi_968,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10x_xi_972,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_992_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_992_inst_req_0;
      type_cast_992_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_992_inst_req_1;
      type_cast_992_inst_ack_1<= rack(0);
      type_cast_992_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_992_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr13x_xi_989,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16x_xi_993,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1179_index_1_rename
    process(R_tmp_1178_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp_1178_resized;
      ov(2 downto 0) := iv;
      R_tmp_1178_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1179_index_1_resize
    process(tmp_1174) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp_1174;
      ov := iv(2 downto 0);
      R_tmp_1178_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1179_root_address_inst
    process(array_obj_ref_1179_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1179_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_1179_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_764_index_1_rename
    process(R_indvar81_763_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar81_763_resized;
      ov(13 downto 0) := iv;
      R_indvar81_763_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_764_index_1_resize
    process(indvar81_752) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar81_752;
      ov := iv(13 downto 0);
      R_indvar81_763_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_764_root_address_inst
    process(array_obj_ref_764_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_764_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_764_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_935_index_1_rename
    process(R_ix_x0x_xlcssa_934_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_934_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_934_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_935_index_1_resize
    process(ix_x0x_xlcssa_900) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_900;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_934_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_935_root_address_inst
    process(array_obj_ref_935_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_935_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_935_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1002_addr_0
    process(ptr_deref_1002_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1002_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1002_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1002_base_resize
    process(arrayidx17x_xi_1000) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx17x_xi_1000;
      ov := iv(2 downto 0);
      ptr_deref_1002_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1002_gather_scatter
    process(conv16x_xi_993) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv16x_xi_993;
      ov(7 downto 0) := iv;
      ptr_deref_1002_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1002_root_address_inst
    process(ptr_deref_1002_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1002_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1002_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1023_addr_0
    process(ptr_deref_1023_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1023_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1023_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1023_base_resize
    process(arrayidx23x_xi_1021) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx23x_xi_1021;
      ov := iv(2 downto 0);
      ptr_deref_1023_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1023_gather_scatter
    process(conv22x_xi_1014) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv22x_xi_1014;
      ov(7 downto 0) := iv;
      ptr_deref_1023_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1023_root_address_inst
    process(ptr_deref_1023_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1023_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1023_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_addr_0
    process(ptr_deref_1044_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1044_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1044_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_base_resize
    process(arrayidx29x_xi_1042) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx29x_xi_1042;
      ov := iv(2 downto 0);
      ptr_deref_1044_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_gather_scatter
    process(conv28x_xi_1035) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv28x_xi_1035;
      ov(7 downto 0) := iv;
      ptr_deref_1044_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_root_address_inst
    process(ptr_deref_1044_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1044_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1044_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1065_addr_0
    process(ptr_deref_1065_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1065_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1065_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1065_base_resize
    process(arrayidx35x_xi_1063) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx35x_xi_1063;
      ov := iv(2 downto 0);
      ptr_deref_1065_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1065_gather_scatter
    process(conv34x_xi_1056) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv34x_xi_1056;
      ov(7 downto 0) := iv;
      ptr_deref_1065_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1065_root_address_inst
    process(ptr_deref_1065_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1065_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1065_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1086_addr_0
    process(ptr_deref_1086_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1086_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1086_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1086_base_resize
    process(arrayidx41x_xi_1084) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx41x_xi_1084;
      ov := iv(2 downto 0);
      ptr_deref_1086_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1086_gather_scatter
    process(conv40x_xi_1077) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv40x_xi_1077;
      ov(7 downto 0) := iv;
      ptr_deref_1086_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1086_root_address_inst
    process(ptr_deref_1086_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1086_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1086_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1183_addr_0
    process(ptr_deref_1183_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1183_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1183_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1183_base_resize
    process(arrayidx49x_xphix_xtransx_xinsertx_xi_1180) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx49x_xphix_xtransx_xinsertx_xi_1180;
      ov := iv(2 downto 0);
      ptr_deref_1183_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1183_gather_scatter
    process(ptr_deref_1183_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1183_data_0;
      ov(7 downto 0) := iv;
      tmp50x_xprex_xi_1184 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1183_root_address_inst
    process(ptr_deref_1183_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1183_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1183_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_769_addr_0
    process(ptr_deref_769_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_769_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_769_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_769_base_resize
    process(arrayidx_766) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_766;
      ov := iv(13 downto 0);
      ptr_deref_769_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_769_gather_scatter
    process(ptr_deref_769_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_769_data_0;
      ov(63 downto 0) := iv;
      tmp4_770 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_769_root_address_inst
    process(ptr_deref_769_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_769_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_769_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_940_addr_0
    process(ptr_deref_940_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_940_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_940_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_940_base_resize
    process(arrayidxx_xi_937) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidxx_xi_937;
      ov := iv(13 downto 0);
      ptr_deref_940_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_940_gather_scatter
    process(ptr_deref_940_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_940_data_0;
      ov(63 downto 0) := iv;
      tmp1x_xi_941 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_940_root_address_inst
    process(ptr_deref_940_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_940_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_940_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_960_addr_0
    process(ptr_deref_960_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_960_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_960_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_960_base_resize
    process(arrayidx5x_xi_958) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx5x_xi_958;
      ov := iv(2 downto 0);
      ptr_deref_960_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_960_gather_scatter
    process(convx_xi_951) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := convx_xi_951;
      ov(7 downto 0) := iv;
      ptr_deref_960_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_960_root_address_inst
    process(ptr_deref_960_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_960_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_960_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_981_addr_0
    process(ptr_deref_981_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_981_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_981_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_981_base_resize
    process(arrayidx11x_xi_979) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx11x_xi_979;
      ov := iv(2 downto 0);
      ptr_deref_981_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_981_gather_scatter
    process(conv10x_xi_972) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv10x_xi_972;
      ov(7 downto 0) := iv;
      ptr_deref_981_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_981_root_address_inst
    process(ptr_deref_981_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_981_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_981_root_address <= ov(2 downto 0);
      --
    end process;
    if_stmt_1095_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp53x_xi_1094;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1095_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1095_branch_req_0,
          ack0 => if_stmt_1095_branch_ack_0,
          ack1 => if_stmt_1095_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1146_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcondx_xi73_1145;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1146_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1146_branch_req_0,
          ack0 => if_stmt_1146_branch_ack_0,
          ack1 => if_stmt_1146_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1193_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_1192;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1193_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1193_branch_req_0,
          ack0 => if_stmt_1193_branch_ack_0,
          ack1 => if_stmt_1193_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_702_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp76_701;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_702_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_702_branch_req_0,
          ack0 => if_stmt_702_branch_ack_0,
          ack1 => if_stmt_702_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_880_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_879;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_880_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_880_branch_req_0,
          ack0 => if_stmt_880_branch_ack_0,
          ack1 => if_stmt_880_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_920_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_919;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_920_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_920_branch_req_0,
          ack0 => if_stmt_920_branch_ack_0,
          ack1 => if_stmt_920_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_738_inst
    process(umax6_733) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(umax6_733, type_cast_737_wire_constant, tmp_var);
      tmp7_739 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1116_inst
    process(tmpx_xi_1105) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmpx_xi_1105, type_cast_1115_wire_constant, tmp_var);
      tmpx_xopx_xi_1117 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1128_inst
    process(iNsTr_30_1123) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_30_1123, type_cast_1127_wire_constant, tmp_var);
      xx_xopx_xi_1129 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1157_inst
    process(tmp58x_xi_1136) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp58x_xi_1136, type_cast_1156_wire_constant, tmp_var);
      tmp2_1158 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1173_inst
    process(indvar1_1161) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar1_1161, type_cast_1172_wire_constant, tmp_var);
      tmp_1174 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1204_inst
    process(indvar1_1161) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar1_1161, type_cast_1203_wire_constant, tmp_var);
      indvarx_xnext_1205 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_748_inst
    process(tmp8_743) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp8_743, type_cast_747_wire_constant, tmp_var);
      tmp9_749 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_873_inst
    process(indvar81_752) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar81_752, type_cast_872_wire_constant, tmp_var);
      indvarx_xnext82_874 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_912_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(size_buffer, type_cast_911_wire_constant, tmp_var);
      and68_913 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1122_inst
    process(tmpx_xopx_xi_1117) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(tmpx_xopx_xi_1117, type_cast_1121_wire_constant, tmp_var);
      iNsTr_30_1123 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_918_inst
    process(and68_913) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and68_913, type_cast_917_wire_constant, tmp_var);
      tobool_919 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1144_inst
    process(tmp58x_xi_1136) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tmp58x_xi_1136, type_cast_1143_wire_constant, tmp_var);
      exitcondx_xi73_1145 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1191_inst
    process(indvar1_1161, tmp2_1158) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvar1_1161, tmp2_1158, tmp_var);
      exitcond3_1192 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_878_inst
    process(indvarx_xnext82_874, tmp9_749) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext82_874, tmp9_749, tmp_var);
      exitcond_879 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1093_inst
    process(conv72_930) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv72_930, type_cast_1092_wire_constant, tmp_var);
      cmp53x_xi_1094 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_713_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(size_buffer, type_cast_712_wire_constant, tmp_var);
      shr_714 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1009_inst
    process(tmp1x_xi_941) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_941, type_cast_1008_wire_constant, tmp_var);
      shr19x_xi_1010 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1030_inst
    process(tmp1x_xi_941) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_941, type_cast_1029_wire_constant, tmp_var);
      shr25x_xi_1031 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1051_inst
    process(tmp1x_xi_941) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_941, type_cast_1050_wire_constant, tmp_var);
      shr31x_xi_1052 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1072_inst
    process(tmp1x_xi_941) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_941, type_cast_1071_wire_constant, tmp_var);
      shr37x_xi_1073 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_779_inst
    process(tmp4_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_770, type_cast_778_wire_constant, tmp_var);
      shr9_780 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_789_inst
    process(tmp4_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_770, type_cast_788_wire_constant, tmp_var);
      shr15_790 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_799_inst
    process(tmp4_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_770, type_cast_798_wire_constant, tmp_var);
      shr21_800 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_809_inst
    process(tmp4_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_770, type_cast_808_wire_constant, tmp_var);
      shr27_810 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_819_inst
    process(tmp4_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_770, type_cast_818_wire_constant, tmp_var);
      shr33_820 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_829_inst
    process(tmp4_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_770, type_cast_828_wire_constant, tmp_var);
      shr39_830 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_839_inst
    process(tmp4_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_770, type_cast_838_wire_constant, tmp_var);
      shr45_840 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_946_inst
    process(tmp1x_xi_941) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_941, type_cast_945_wire_constant, tmp_var);
      shrx_xi_947 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_967_inst
    process(tmp1x_xi_941) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_941, type_cast_966_wire_constant, tmp_var);
      shr7x_xi_968 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_988_inst
    process(tmp1x_xi_941) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_941, type_cast_987_wire_constant, tmp_var);
      shr13x_xi_989 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_700_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(size_buffer, type_cast_699_wire_constant, tmp_var);
      cmp76_701 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_719_inst
    process(shr_714) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_714, type_cast_718_wire_constant, tmp_var);
      tmp80_720 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_725_inst
    process(shr_714) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_714, type_cast_724_wire_constant, tmp_var);
      tmp5_726 <= tmp_var; --
    end process;
    -- binary operator UGT_u8_u1_1110_inst
    process(conv72_930) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv72_930, type_cast_1109_wire_constant, tmp_var);
      tmp55x_xi_1111 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_1179_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_tmp_1178_scaled;
      array_obj_ref_1179_final_offset <= data_out(2 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1179_index_offset_req_0;
      array_obj_ref_1179_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1179_index_offset_req_1;
      array_obj_ref_1179_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_764_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar81_763_scaled;
      array_obj_ref_764_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_764_index_offset_req_0;
      array_obj_ref_764_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_764_index_offset_req_1;
      array_obj_ref_764_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_935_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_934_scaled;
      array_obj_ref_935_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_935_index_offset_req_0;
      array_obj_ref_935_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_935_index_offset_req_1;
      array_obj_ref_935_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared load operator group (0) : ptr_deref_1183_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1183_load_0_req_0;
      ptr_deref_1183_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1183_load_0_req_1;
      ptr_deref_1183_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1183_word_address_0;
      ptr_deref_1183_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 3,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(2 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(7 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_940_load_0 ptr_deref_769_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_940_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_769_load_0_req_0;
      ptr_deref_940_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_769_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_940_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_769_load_0_req_1;
      ptr_deref_940_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_769_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_940_word_address_0 & ptr_deref_769_word_address_0;
      ptr_deref_940_data_0 <= data_out(127 downto 64);
      ptr_deref_769_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : ptr_deref_1044_store_0 ptr_deref_960_store_0 ptr_deref_1023_store_0 ptr_deref_1002_store_0 ptr_deref_981_store_0 ptr_deref_1086_store_0 ptr_deref_1065_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(55 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= ptr_deref_1044_store_0_req_0;
      reqL_unguarded(5) <= ptr_deref_960_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1023_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_1002_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_981_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1086_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1065_store_0_req_0;
      ptr_deref_1044_store_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_960_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1023_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_1002_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_981_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1086_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1065_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= ptr_deref_1044_store_0_req_1;
      reqR_unguarded(5) <= ptr_deref_960_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1023_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_1002_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_981_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1086_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1065_store_0_req_1;
      ptr_deref_1044_store_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_960_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1023_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_1002_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_981_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1086_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1065_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_6: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1044_word_address_0 & ptr_deref_960_word_address_0 & ptr_deref_1023_word_address_0 & ptr_deref_1002_word_address_0 & ptr_deref_981_word_address_0 & ptr_deref_1086_word_address_0 & ptr_deref_1065_word_address_0;
      data_in <= ptr_deref_1044_data_0 & ptr_deref_960_data_0 & ptr_deref_1023_data_0 & ptr_deref_1002_data_0 & ptr_deref_981_data_0 & ptr_deref_1086_data_0 & ptr_deref_1065_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 3,
        data_width => 8,
        num_reqs => 7,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(2 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 7,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_860_inst WPIPE_maxpool_output_pipe_866_inst WPIPE_maxpool_output_pipe_857_inst WPIPE_maxpool_output_pipe_854_inst WPIPE_maxpool_output_pipe_1137_inst WPIPE_maxpool_output_pipe_863_inst WPIPE_maxpool_output_pipe_851_inst WPIPE_maxpool_output_pipe_848_inst WPIPE_maxpool_output_pipe_845_inst WPIPE_maxpool_output_pipe_1185_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal sample_req, sample_ack : BooleanArray( 9 downto 0);
      signal update_req, update_ack : BooleanArray( 9 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 9 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 9 downto 0);
      signal guard_vector : std_logic_vector( 9 downto 0);
      constant inBUFs : IntegerArray(9 downto 0) := (9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(9 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false);
      constant guardBuffering: IntegerArray(9 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2);
      -- 
    begin -- 
      sample_req_unguarded(9) <= WPIPE_maxpool_output_pipe_860_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_maxpool_output_pipe_866_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_857_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_854_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1137_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_863_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_851_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_848_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_845_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1185_inst_req_0;
      WPIPE_maxpool_output_pipe_860_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_866_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_857_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_854_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1137_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_863_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_851_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_848_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_845_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1185_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(9) <= WPIPE_maxpool_output_pipe_860_inst_req_1;
      update_req_unguarded(8) <= WPIPE_maxpool_output_pipe_866_inst_req_1;
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_857_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_854_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1137_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_863_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_851_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_848_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_845_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1185_inst_req_1;
      WPIPE_maxpool_output_pipe_860_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_866_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_857_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_854_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1137_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_863_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_851_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_848_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_845_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1185_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      data_in <= conv18_794 & conv_774 & conv24_804 & conv30_814 & conv40x_xi_1077 & conv12_784 & conv36_824 & conv42_834 & conv48_844 & tmp50x_xprex_xi_1184;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 10, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 10, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 1,
      addr_width => 3,
      data_width => 8,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 3,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end sendB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendModule is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    output_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
    output_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
    output_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendModule;
architecture sendModule_arch of sendModule is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendModule_CP_7983_start: Boolean;
  signal sendModule_CP_7983_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_3303_load_0_ack_0 : boolean;
  signal ptr_deref_3303_load_0_req_0 : boolean;
  signal slice_3310_inst_req_0 : boolean;
  signal slice_3310_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3306_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3306_inst_ack_0 : boolean;
  signal EQ_u3_u1_3517_inst_ack_0 : boolean;
  signal ptr_deref_3303_load_0_ack_1 : boolean;
  signal ptr_deref_3303_load_0_req_1 : boolean;
  signal slice_3314_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3306_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3306_inst_ack_1 : boolean;
  signal slice_3310_inst_req_1 : boolean;
  signal slice_3310_inst_ack_1 : boolean;
  signal slice_3314_inst_req_1 : boolean;
  signal slice_3314_inst_ack_1 : boolean;
  signal W_output_data2_3338_delayed_13_0_3519_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3147_inst_req_0 : boolean;
  signal EQ_u3_u1_3545_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3147_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3147_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3147_inst_ack_1 : boolean;
  signal EQ_u3_u1_3545_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_3631_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3150_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3150_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3150_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3150_inst_ack_1 : boolean;
  signal EQ_u3_u1_3545_inst_req_1 : boolean;
  signal EQ_u3_u1_3545_inst_ack_1 : boolean;
  signal RPIPE_output_pipe_3153_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3153_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3153_inst_req_1 : boolean;
  signal W_output_data2_3378_delayed_13_0_3589_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3153_inst_ack_1 : boolean;
  signal W_fetch_addr2_3408_delayed_8_0_3633_inst_ack_1 : boolean;
  signal do_while_stmt_3161_branch_req_0 : boolean;
  signal W_output_data2_3338_delayed_13_0_3519_inst_ack_0 : boolean;
  signal W_output_data2_3330_delayed_13_0_3505_inst_req_0 : boolean;
  signal EQ_u3_u1_3531_inst_ack_0 : boolean;
  signal phi_stmt_3163_req_1 : boolean;
  signal W_output_data2_3330_delayed_13_0_3505_inst_ack_0 : boolean;
  signal EQ_u3_u1_3573_inst_req_1 : boolean;
  signal W_output_data2_3354_delayed_13_0_3547_inst_req_0 : boolean;
  signal phi_stmt_3163_req_0 : boolean;
  signal phi_stmt_3163_ack_0 : boolean;
  signal W_output_data2_3354_delayed_13_0_3547_inst_ack_0 : boolean;
  signal EQ_u3_u1_3531_inst_req_1 : boolean;
  signal W_fetch_addr1_3390_delayed_8_0_3612_inst_req_0 : boolean;
  signal W_fetch_addr1_3390_delayed_8_0_3612_inst_ack_0 : boolean;
  signal W_output_data2_3354_delayed_13_0_3547_inst_req_1 : boolean;
  signal n_address1_3262_3167_buf_req_0 : boolean;
  signal n_address1_3262_3167_buf_ack_0 : boolean;
  signal W_output_data2_3338_delayed_13_0_3519_inst_req_1 : boolean;
  signal W_output_data2_3354_delayed_13_0_3547_inst_ack_1 : boolean;
  signal n_address1_3262_3167_buf_req_1 : boolean;
  signal W_output_data2_3378_delayed_13_0_3589_inst_ack_1 : boolean;
  signal n_address1_3262_3167_buf_ack_1 : boolean;
  signal W_output_data2_3338_delayed_13_0_3519_inst_ack_1 : boolean;
  signal phi_stmt_3168_req_1 : boolean;
  signal phi_stmt_3168_req_0 : boolean;
  signal EQ_u3_u1_3531_inst_ack_1 : boolean;
  signal W_fetch_addr1_3390_delayed_8_0_3612_inst_req_1 : boolean;
  signal phi_stmt_3168_ack_0 : boolean;
  signal W_output_data2_3330_delayed_13_0_3505_inst_req_1 : boolean;
  signal W_fetch_addr1_3390_delayed_8_0_3612_inst_ack_1 : boolean;
  signal W_output_data2_3330_delayed_13_0_3505_inst_ack_1 : boolean;
  signal type_cast_3171_inst_req_0 : boolean;
  signal type_cast_3171_inst_ack_0 : boolean;
  signal type_cast_3171_inst_req_1 : boolean;
  signal type_cast_3171_inst_ack_1 : boolean;
  signal n_address2_3276_3172_buf_req_0 : boolean;
  signal n_address2_3276_3172_buf_ack_0 : boolean;
  signal EQ_u3_u1_3573_inst_ack_1 : boolean;
  signal EQ_u3_u1_3559_inst_req_0 : boolean;
  signal n_address2_3276_3172_buf_req_1 : boolean;
  signal EQ_u3_u1_3559_inst_ack_0 : boolean;
  signal n_address2_3276_3172_buf_ack_1 : boolean;
  signal EQ_u3_u1_3559_inst_req_1 : boolean;
  signal EQ_u3_u1_3559_inst_ack_1 : boolean;
  signal phi_stmt_3173_req_1 : boolean;
  signal phi_stmt_3173_req_0 : boolean;
  signal phi_stmt_3173_ack_0 : boolean;
  signal W_output_data2_3362_delayed_13_0_3561_inst_req_0 : boolean;
  signal n_chl_3232_3177_buf_req_0 : boolean;
  signal n_chl_3232_3177_buf_ack_0 : boolean;
  signal CONCAT_u32_u64_3631_inst_req_1 : boolean;
  signal n_chl_3232_3177_buf_req_1 : boolean;
  signal n_chl_3232_3177_buf_ack_1 : boolean;
  signal W_output_data2_3362_delayed_13_0_3561_inst_ack_0 : boolean;
  signal EQ_u3_u1_3517_inst_req_1 : boolean;
  signal W_output_data2_3362_delayed_13_0_3561_inst_req_1 : boolean;
  signal phi_stmt_3178_req_1 : boolean;
  signal EQ_u3_u1_3601_inst_req_0 : boolean;
  signal phi_stmt_3178_req_0 : boolean;
  signal slice_3314_inst_ack_0 : boolean;
  signal W_output_data2_3362_delayed_13_0_3561_inst_ack_1 : boolean;
  signal phi_stmt_3178_ack_0 : boolean;
  signal CONCAT_u32_u64_3652_inst_req_0 : boolean;
  signal CONCAT_u32_u64_3631_inst_req_0 : boolean;
  signal n_col_3213_3182_buf_req_0 : boolean;
  signal EQ_u3_u1_3601_inst_ack_0 : boolean;
  signal n_col_3213_3182_buf_ack_0 : boolean;
  signal n_col_3213_3182_buf_req_1 : boolean;
  signal n_col_3213_3182_buf_ack_1 : boolean;
  signal EQ_u3_u1_3531_inst_req_0 : boolean;
  signal phi_stmt_3183_req_1 : boolean;
  signal phi_stmt_3183_req_0 : boolean;
  signal phi_stmt_3183_ack_0 : boolean;
  signal n_row_3224_3187_buf_req_0 : boolean;
  signal n_row_3224_3187_buf_ack_0 : boolean;
  signal n_row_3224_3187_buf_req_1 : boolean;
  signal n_row_3224_3187_buf_ack_1 : boolean;
  signal SUB_u16_u16_3197_inst_req_0 : boolean;
  signal SUB_u16_u16_3197_inst_ack_0 : boolean;
  signal SUB_u16_u16_3197_inst_req_1 : boolean;
  signal SUB_u16_u16_3197_inst_ack_1 : boolean;
  signal type_cast_3235_inst_req_0 : boolean;
  signal type_cast_3235_inst_ack_0 : boolean;
  signal type_cast_3235_inst_req_1 : boolean;
  signal type_cast_3235_inst_ack_1 : boolean;
  signal type_cast_3244_inst_req_0 : boolean;
  signal type_cast_3244_inst_ack_0 : boolean;
  signal type_cast_3244_inst_req_1 : boolean;
  signal type_cast_3244_inst_ack_1 : boolean;
  signal array_obj_ref_3284_index_offset_req_0 : boolean;
  signal array_obj_ref_3284_index_offset_ack_0 : boolean;
  signal array_obj_ref_3284_index_offset_req_1 : boolean;
  signal array_obj_ref_3284_index_offset_ack_1 : boolean;
  signal addr_of_3285_final_reg_req_0 : boolean;
  signal addr_of_3285_final_reg_ack_0 : boolean;
  signal addr_of_3285_final_reg_req_1 : boolean;
  signal addr_of_3285_final_reg_ack_1 : boolean;
  signal array_obj_ref_3294_index_offset_req_0 : boolean;
  signal array_obj_ref_3294_index_offset_ack_0 : boolean;
  signal array_obj_ref_3294_index_offset_req_1 : boolean;
  signal array_obj_ref_3294_index_offset_ack_1 : boolean;
  signal addr_of_3295_final_reg_req_0 : boolean;
  signal addr_of_3295_final_reg_ack_0 : boolean;
  signal addr_of_3295_final_reg_req_1 : boolean;
  signal addr_of_3295_final_reg_ack_1 : boolean;
  signal ptr_deref_3299_load_0_req_0 : boolean;
  signal ptr_deref_3299_load_0_ack_0 : boolean;
  signal ptr_deref_3299_load_0_req_1 : boolean;
  signal ptr_deref_3299_load_0_ack_1 : boolean;
  signal slice_3318_inst_req_0 : boolean;
  signal slice_3318_inst_ack_0 : boolean;
  signal slice_3318_inst_req_1 : boolean;
  signal slice_3318_inst_ack_1 : boolean;
  signal slice_3322_inst_req_0 : boolean;
  signal slice_3322_inst_ack_0 : boolean;
  signal slice_3322_inst_req_1 : boolean;
  signal slice_3322_inst_ack_1 : boolean;
  signal slice_3326_inst_req_0 : boolean;
  signal slice_3326_inst_ack_0 : boolean;
  signal slice_3326_inst_req_1 : boolean;
  signal slice_3326_inst_ack_1 : boolean;
  signal slice_3330_inst_req_0 : boolean;
  signal slice_3330_inst_ack_0 : boolean;
  signal slice_3330_inst_req_1 : boolean;
  signal slice_3330_inst_ack_1 : boolean;
  signal slice_3334_inst_req_0 : boolean;
  signal slice_3334_inst_ack_0 : boolean;
  signal slice_3334_inst_req_1 : boolean;
  signal slice_3334_inst_ack_1 : boolean;
  signal slice_3338_inst_req_0 : boolean;
  signal slice_3338_inst_ack_0 : boolean;
  signal slice_3338_inst_req_1 : boolean;
  signal slice_3338_inst_ack_1 : boolean;
  signal slice_3342_inst_req_0 : boolean;
  signal slice_3342_inst_ack_0 : boolean;
  signal slice_3342_inst_req_1 : boolean;
  signal slice_3342_inst_ack_1 : boolean;
  signal slice_3346_inst_req_0 : boolean;
  signal slice_3346_inst_ack_0 : boolean;
  signal slice_3346_inst_req_1 : boolean;
  signal slice_3346_inst_ack_1 : boolean;
  signal slice_3350_inst_req_0 : boolean;
  signal slice_3350_inst_ack_0 : boolean;
  signal slice_3350_inst_req_1 : boolean;
  signal slice_3350_inst_ack_1 : boolean;
  signal slice_3354_inst_req_0 : boolean;
  signal slice_3354_inst_ack_0 : boolean;
  signal slice_3354_inst_req_1 : boolean;
  signal slice_3354_inst_ack_1 : boolean;
  signal slice_3358_inst_req_0 : boolean;
  signal slice_3358_inst_ack_0 : boolean;
  signal slice_3358_inst_req_1 : boolean;
  signal slice_3358_inst_ack_1 : boolean;
  signal slice_3362_inst_req_0 : boolean;
  signal slice_3362_inst_ack_0 : boolean;
  signal slice_3362_inst_req_1 : boolean;
  signal slice_3362_inst_ack_1 : boolean;
  signal slice_3366_inst_req_0 : boolean;
  signal slice_3366_inst_ack_0 : boolean;
  signal slice_3366_inst_req_1 : boolean;
  signal slice_3366_inst_ack_1 : boolean;
  signal slice_3370_inst_req_0 : boolean;
  signal slice_3370_inst_ack_0 : boolean;
  signal slice_3370_inst_req_1 : boolean;
  signal slice_3370_inst_ack_1 : boolean;
  signal slice_3374_inst_req_0 : boolean;
  signal slice_3374_inst_ack_0 : boolean;
  signal slice_3374_inst_req_1 : boolean;
  signal slice_3374_inst_ack_1 : boolean;
  signal slice_3378_inst_req_0 : boolean;
  signal slice_3378_inst_ack_0 : boolean;
  signal slice_3378_inst_req_1 : boolean;
  signal slice_3378_inst_ack_1 : boolean;
  signal EQ_u3_u1_3391_inst_req_0 : boolean;
  signal EQ_u3_u1_3391_inst_ack_0 : boolean;
  signal W_fetch_addr2_3408_delayed_8_0_3633_inst_req_1 : boolean;
  signal EQ_u3_u1_3391_inst_req_1 : boolean;
  signal EQ_u3_u1_3391_inst_ack_1 : boolean;
  signal W_output_data1_3266_delayed_13_0_3393_inst_req_0 : boolean;
  signal W_output_data2_3378_delayed_13_0_3589_inst_ack_0 : boolean;
  signal W_output_data1_3266_delayed_13_0_3393_inst_ack_0 : boolean;
  signal W_output_data1_3266_delayed_13_0_3393_inst_req_1 : boolean;
  signal W_output_data2_3378_delayed_13_0_3589_inst_req_0 : boolean;
  signal W_output_data1_3266_delayed_13_0_3393_inst_ack_1 : boolean;
  signal W_fetch_addr2_3408_delayed_8_0_3633_inst_ack_0 : boolean;
  signal W_fetch_addr2_3408_delayed_8_0_3633_inst_req_0 : boolean;
  signal EQ_u3_u1_3405_inst_req_0 : boolean;
  signal EQ_u3_u1_3405_inst_ack_0 : boolean;
  signal EQ_u3_u1_3573_inst_ack_0 : boolean;
  signal EQ_u3_u1_3405_inst_req_1 : boolean;
  signal EQ_u3_u1_3405_inst_ack_1 : boolean;
  signal EQ_u3_u1_3517_inst_req_0 : boolean;
  signal W_output_data2_3386_delayed_13_0_3603_inst_ack_1 : boolean;
  signal W_output_data1_3274_delayed_13_0_3407_inst_req_0 : boolean;
  signal W_output_data1_3274_delayed_13_0_3407_inst_ack_0 : boolean;
  signal W_output_data1_3274_delayed_13_0_3407_inst_req_1 : boolean;
  signal W_output_data1_3274_delayed_13_0_3407_inst_ack_1 : boolean;
  signal W_output_data2_3386_delayed_13_0_3603_inst_req_1 : boolean;
  signal EQ_u3_u1_3419_inst_req_0 : boolean;
  signal EQ_u3_u1_3419_inst_ack_0 : boolean;
  signal EQ_u3_u1_3419_inst_req_1 : boolean;
  signal EQ_u3_u1_3587_inst_ack_1 : boolean;
  signal EQ_u3_u1_3419_inst_ack_1 : boolean;
  signal ptr_deref_3616_store_0_ack_1 : boolean;
  signal W_output_data1_3282_delayed_13_0_3421_inst_req_0 : boolean;
  signal EQ_u3_u1_3587_inst_req_1 : boolean;
  signal W_output_data1_3282_delayed_13_0_3421_inst_ack_0 : boolean;
  signal ptr_deref_3616_store_0_req_1 : boolean;
  signal W_output_data1_3282_delayed_13_0_3421_inst_req_1 : boolean;
  signal W_output_data1_3282_delayed_13_0_3421_inst_ack_1 : boolean;
  signal W_output_data2_3386_delayed_13_0_3603_inst_ack_0 : boolean;
  signal W_output_data2_3346_delayed_13_0_3533_inst_ack_1 : boolean;
  signal EQ_u3_u1_3433_inst_req_0 : boolean;
  signal EQ_u3_u1_3587_inst_ack_0 : boolean;
  signal EQ_u3_u1_3433_inst_ack_0 : boolean;
  signal EQ_u3_u1_3573_inst_req_0 : boolean;
  signal EQ_u3_u1_3433_inst_req_1 : boolean;
  signal EQ_u3_u1_3587_inst_req_0 : boolean;
  signal EQ_u3_u1_3433_inst_ack_1 : boolean;
  signal W_output_data2_3386_delayed_13_0_3603_inst_req_0 : boolean;
  signal W_output_data2_3346_delayed_13_0_3533_inst_req_1 : boolean;
  signal W_output_data1_3290_delayed_13_0_3435_inst_req_0 : boolean;
  signal W_output_data1_3290_delayed_13_0_3435_inst_ack_0 : boolean;
  signal W_output_data1_3290_delayed_13_0_3435_inst_req_1 : boolean;
  signal W_output_data1_3290_delayed_13_0_3435_inst_ack_1 : boolean;
  signal ptr_deref_3616_store_0_ack_0 : boolean;
  signal EQ_u3_u1_3447_inst_req_0 : boolean;
  signal EQ_u3_u1_3447_inst_ack_0 : boolean;
  signal ptr_deref_3616_store_0_req_0 : boolean;
  signal EQ_u3_u1_3447_inst_req_1 : boolean;
  signal EQ_u3_u1_3447_inst_ack_1 : boolean;
  signal W_output_data1_3298_delayed_13_0_3449_inst_req_0 : boolean;
  signal W_output_data1_3298_delayed_13_0_3449_inst_ack_0 : boolean;
  signal W_output_data1_3298_delayed_13_0_3449_inst_req_1 : boolean;
  signal W_output_data2_3370_delayed_13_0_3575_inst_ack_1 : boolean;
  signal W_output_data1_3298_delayed_13_0_3449_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_3652_inst_ack_1 : boolean;
  signal EQ_u3_u1_3503_inst_ack_1 : boolean;
  signal W_output_data2_3370_delayed_13_0_3575_inst_req_1 : boolean;
  signal EQ_u3_u1_3461_inst_req_0 : boolean;
  signal EQ_u3_u1_3461_inst_ack_0 : boolean;
  signal EQ_u3_u1_3461_inst_req_1 : boolean;
  signal EQ_u3_u1_3461_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_3652_inst_req_1 : boolean;
  signal W_output_data2_3346_delayed_13_0_3533_inst_ack_0 : boolean;
  signal W_output_data1_3306_delayed_13_0_3463_inst_req_0 : boolean;
  signal W_output_data2_3370_delayed_13_0_3575_inst_ack_0 : boolean;
  signal W_output_data1_3306_delayed_13_0_3463_inst_ack_0 : boolean;
  signal W_output_data1_3306_delayed_13_0_3463_inst_req_1 : boolean;
  signal W_output_data2_3370_delayed_13_0_3575_inst_req_0 : boolean;
  signal W_output_data1_3306_delayed_13_0_3463_inst_ack_1 : boolean;
  signal EQ_u3_u1_3601_inst_ack_1 : boolean;
  signal W_output_data2_3346_delayed_13_0_3533_inst_req_0 : boolean;
  signal EQ_u3_u1_3503_inst_req_1 : boolean;
  signal EQ_u3_u1_3475_inst_req_0 : boolean;
  signal EQ_u3_u1_3475_inst_ack_0 : boolean;
  signal EQ_u3_u1_3475_inst_req_1 : boolean;
  signal EQ_u3_u1_3475_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_3652_inst_ack_0 : boolean;
  signal EQ_u3_u1_3601_inst_req_1 : boolean;
  signal CONCAT_u32_u64_3631_inst_ack_1 : boolean;
  signal W_output_data1_3314_delayed_13_0_3477_inst_req_0 : boolean;
  signal W_output_data1_3314_delayed_13_0_3477_inst_ack_0 : boolean;
  signal W_output_data1_3314_delayed_13_0_3477_inst_req_1 : boolean;
  signal W_output_data1_3314_delayed_13_0_3477_inst_ack_1 : boolean;
  signal EQ_u3_u1_3517_inst_ack_1 : boolean;
  signal EQ_u3_u1_3489_inst_req_0 : boolean;
  signal EQ_u3_u1_3489_inst_ack_0 : boolean;
  signal EQ_u3_u1_3489_inst_req_1 : boolean;
  signal EQ_u3_u1_3489_inst_ack_1 : boolean;
  signal W_output_data1_3322_delayed_13_0_3491_inst_req_0 : boolean;
  signal W_output_data1_3322_delayed_13_0_3491_inst_ack_0 : boolean;
  signal W_output_data1_3322_delayed_13_0_3491_inst_req_1 : boolean;
  signal W_output_data1_3322_delayed_13_0_3491_inst_ack_1 : boolean;
  signal EQ_u3_u1_3503_inst_req_0 : boolean;
  signal EQ_u3_u1_3503_inst_ack_0 : boolean;
  signal ptr_deref_3637_store_0_req_0 : boolean;
  signal ptr_deref_3637_store_0_ack_0 : boolean;
  signal ptr_deref_3637_store_0_req_1 : boolean;
  signal ptr_deref_3637_store_0_ack_1 : boolean;
  signal SUB_u16_u16_3657_inst_req_0 : boolean;
  signal SUB_u16_u16_3657_inst_ack_0 : boolean;
  signal SUB_u16_u16_3657_inst_req_1 : boolean;
  signal SUB_u16_u16_3657_inst_ack_1 : boolean;
  signal do_while_stmt_3161_branch_ack_0 : boolean;
  signal do_while_stmt_3161_branch_ack_1 : boolean;
  signal WPIPE_input_done_pipe_3669_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_3669_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_3669_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_3669_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendModule_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendModule_CP_7983_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendModule_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendModule_CP_7983_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendModule_CP_7983_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendModule_CP_7983_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendModule_CP_7983: Block -- control-path 
    signal sendModule_CP_7983_elements: BooleanArray(391 downto 0);
    -- 
  begin -- 
    sendModule_CP_7983_elements(0) <= sendModule_CP_7983_start;
    sendModule_CP_7983_symbol <= sendModule_CP_7983_elements(391);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_3145/$entry
      -- CP-element group 0: 	 branch_block_stmt_3145/branch_block_stmt_3145__entry__
      -- CP-element group 0: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160__entry__
      -- CP-element group 0: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/$entry
      -- CP-element group 0: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_Sample/rr
      -- 
    rr_8007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(0), ack => RPIPE_output_pipe_3147_inst_req_0); -- 
    -- CP-element group 1:  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	389 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	390 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_3145/do_while_stmt_3161__exit__
      -- CP-element group 1: 	 branch_block_stmt_3145/assign_stmt_3671__entry__
      -- CP-element group 1: 	 branch_block_stmt_3145/assign_stmt_3671/$entry
      -- CP-element group 1: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_Sample/req
      -- 
    req_9434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(1), ack => WPIPE_input_done_pipe_3669_inst_req_0); -- 
    sendModule_CP_7983_elements(1) <= sendModule_CP_7983_elements(389);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_update_start_
      -- CP-element group 2: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_Update/cr
      -- 
    ra_8008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3147_inst_ack_0, ack => sendModule_CP_7983_elements(2)); -- 
    cr_8012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(2), ack => RPIPE_output_pipe_3147_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3147_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_Sample/rr
      -- 
    ca_8013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3147_inst_ack_1, ack => sendModule_CP_7983_elements(3)); -- 
    rr_8021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(3), ack => RPIPE_output_pipe_3150_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_update_start_
      -- CP-element group 4: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_Update/cr
      -- 
    ra_8022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3150_inst_ack_0, ack => sendModule_CP_7983_elements(4)); -- 
    cr_8026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(4), ack => RPIPE_output_pipe_3150_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3150_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_Sample/rr
      -- 
    ca_8027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3150_inst_ack_1, ack => sendModule_CP_7983_elements(5)); -- 
    rr_8035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(5), ack => RPIPE_output_pipe_3153_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_update_start_
      -- CP-element group 6: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_Update/cr
      -- 
    ra_8036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3153_inst_ack_0, ack => sendModule_CP_7983_elements(6)); -- 
    cr_8040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(6), ack => RPIPE_output_pipe_3153_inst_req_1); -- 
    -- CP-element group 7:  transition  place  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160__exit__
      -- CP-element group 7: 	 branch_block_stmt_3145/do_while_stmt_3161__entry__
      -- CP-element group 7: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/$exit
      -- CP-element group 7: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_3145/assign_stmt_3148_to_assign_stmt_3160/RPIPE_output_pipe_3153_Update/ca
      -- 
    ca_8041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3153_inst_ack_1, ack => sendModule_CP_7983_elements(7)); -- 
    -- CP-element group 8:  transition  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_3145/do_while_stmt_3161/$entry
      -- CP-element group 8: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161__entry__
      -- 
    sendModule_CP_7983_elements(8) <= sendModule_CP_7983_elements(7);
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	389 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161__exit__
      -- 
    -- Element group sendModule_CP_7983_elements(9) is bound as output of CP function.
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_3145/do_while_stmt_3161/loop_back
      -- 
    -- Element group sendModule_CP_7983_elements(10) is bound as output of CP function.
    -- CP-element group 11:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	387 
    -- CP-element group 11: 	388 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_3145/do_while_stmt_3161/condition_done
      -- CP-element group 11: 	 branch_block_stmt_3145/do_while_stmt_3161/loop_exit/$entry
      -- CP-element group 11: 	 branch_block_stmt_3145/do_while_stmt_3161/loop_taken/$entry
      -- 
    sendModule_CP_7983_elements(11) <= sendModule_CP_7983_elements(16);
    -- CP-element group 12:  branch  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	386 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_3145/do_while_stmt_3161/loop_body_done
      -- 
    sendModule_CP_7983_elements(12) <= sendModule_CP_7983_elements(386);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	25 
    -- CP-element group 13: 	44 
    -- CP-element group 13: 	65 
    -- CP-element group 13: 	84 
    -- CP-element group 13: 	103 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/back_edge_to_loop_body
      -- 
    sendModule_CP_7983_elements(13) <= sendModule_CP_7983_elements(10);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	27 
    -- CP-element group 14: 	46 
    -- CP-element group 14: 	67 
    -- CP-element group 14: 	86 
    -- CP-element group 14: 	105 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/first_time_through_loop_body
      -- 
    sendModule_CP_7983_elements(14) <= sendModule_CP_7983_elements(8);
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	39 
    -- CP-element group 15: 	59 
    -- CP-element group 15: 	60 
    -- CP-element group 15: 	78 
    -- CP-element group 15: 	79 
    -- CP-element group 15: 	97 
    -- CP-element group 15: 	98 
    -- CP-element group 15: 	137 
    -- CP-element group 15: 	378 
    -- CP-element group 15: 	382 
    -- CP-element group 15: 	150 
    -- CP-element group 15: 	116 
    -- CP-element group 15: 	120 
    -- CP-element group 15: 	124 
    -- CP-element group 15: 	129 
    -- CP-element group 15: 	130 
    -- CP-element group 15: 	136 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/$entry
      -- CP-element group 15: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/loop_body_start
      -- 
    -- Element group sendModule_CP_7983_elements(15) is bound as output of CP function.
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	381 
    -- CP-element group 16: 	382 
    -- CP-element group 16: 	119 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/condition_evaluated
      -- 
    condition_evaluated_8056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_8056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(16), ack => do_while_stmt_3161_branch_req_0); -- 
    sendModule_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(20) & sendModule_CP_7983_elements(381) & sendModule_CP_7983_elements(382) & sendModule_CP_7983_elements(119);
      gj_sendModule_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	21 
    -- CP-element group 17: 	38 
    -- CP-element group 17: 	59 
    -- CP-element group 17: 	78 
    -- CP-element group 17: 	97 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	40 
    -- CP-element group 17: 	61 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	99 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/aggregated_phi_sample_req
      -- CP-element group 17: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_sample_start__ps
      -- 
    sendModule_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(21) & sendModule_CP_7983_elements(38) & sendModule_CP_7983_elements(59) & sendModule_CP_7983_elements(78) & sendModule_CP_7983_elements(97) & sendModule_CP_7983_elements(20);
      gj_sendModule_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	23 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	81 
    -- CP-element group 18: 	100 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	386 
    -- CP-element group 18: 	117 
    -- CP-element group 18: 	121 
    -- CP-element group 18: 	125 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	38 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	78 
    -- CP-element group 18: 	97 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/aggregated_phi_sample_ack
      -- CP-element group 18: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_sample_completed_
      -- 
    sendModule_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(23) & sendModule_CP_7983_elements(41) & sendModule_CP_7983_elements(62) & sendModule_CP_7983_elements(81) & sendModule_CP_7983_elements(100);
      gj_sendModule_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	39 
    -- CP-element group 19: 	60 
    -- CP-element group 19: 	79 
    -- CP-element group 19: 	98 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	63 
    -- CP-element group 19: 	82 
    -- CP-element group 19: 	101 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/aggregated_phi_update_req
      -- CP-element group 19: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_update_start__ps
      -- 
    sendModule_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(22) & sendModule_CP_7983_elements(39) & sendModule_CP_7983_elements(60) & sendModule_CP_7983_elements(79) & sendModule_CP_7983_elements(98);
      gj_sendModule_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	64 
    -- CP-element group 20: 	83 
    -- CP-element group 20: 	102 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/aggregated_phi_update_ack
      -- 
    sendModule_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(24) & sendModule_CP_7983_elements(43) & sendModule_CP_7983_elements(64) & sendModule_CP_7983_elements(83) & sendModule_CP_7983_elements(102);
      gj_sendModule_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: 	119 
    -- CP-element group 21: 	123 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_sample_start_
      -- 
    sendModule_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(18) & sendModule_CP_7983_elements(119) & sendModule_CP_7983_elements(123);
      gj_sendModule_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	268 
    -- CP-element group 22: 	276 
    -- CP-element group 22: 	284 
    -- CP-element group 22: 	252 
    -- CP-element group 22: 	260 
    -- CP-element group 22: 	236 
    -- CP-element group 22: 	244 
    -- CP-element group 22: 	228 
    -- CP-element group 22: 	131 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	19 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_update_start_
      -- 
    sendModule_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(268) & sendModule_CP_7983_elements(276) & sendModule_CP_7983_elements(284) & sendModule_CP_7983_elements(252) & sendModule_CP_7983_elements(260) & sendModule_CP_7983_elements(236) & sendModule_CP_7983_elements(244) & sendModule_CP_7983_elements(228) & sendModule_CP_7983_elements(131);
      gj_sendModule_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	18 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7983_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24: 	274 
    -- CP-element group 24: 	282 
    -- CP-element group 24: 	250 
    -- CP-element group 24: 	258 
    -- CP-element group 24: 	266 
    -- CP-element group 24: 	234 
    -- CP-element group 24: 	242 
    -- CP-element group 24: 	226 
    -- CP-element group 24: 	131 
    -- CP-element group 24:  members (15) 
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_update_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_resized_1
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_scaled_1
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_computed_1
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_resize_1/$entry
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_resize_1/$exit
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_resize_1/index_resize_req
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_resize_1/index_resize_ack
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_scale_1/$entry
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_scale_1/$exit
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_scale_1/scale_rename_req
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_index_scale_1/scale_rename_ack
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_final_index_sum_regn_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_final_index_sum_regn_Sample/req
      -- 
    req_8358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(24), ack => array_obj_ref_3284_index_offset_req_0); -- 
    -- Element group sendModule_CP_7983_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	13 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_loopback_trigger
      -- 
    sendModule_CP_7983_elements(25) <= sendModule_CP_7983_elements(13);
    -- CP-element group 26:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_loopback_sample_req
      -- CP-element group 26: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_loopback_sample_req_ps
      -- 
    phi_stmt_3163_loopback_sample_req_8071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3163_loopback_sample_req_8071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(26), ack => phi_stmt_3163_req_1); -- 
    -- Element group sendModule_CP_7983_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	14 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_entry_trigger
      -- 
    sendModule_CP_7983_elements(27) <= sendModule_CP_7983_elements(14);
    -- CP-element group 28:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_entry_sample_req
      -- CP-element group 28: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_entry_sample_req_ps
      -- 
    phi_stmt_3163_entry_sample_req_8074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3163_entry_sample_req_8074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(28), ack => phi_stmt_3163_req_0); -- 
    -- Element group sendModule_CP_7983_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_phi_mux_ack
      -- CP-element group 29: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3163_phi_mux_ack_ps
      -- 
    phi_stmt_3163_phi_mux_ack_8077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3163_ack_0, ack => sendModule_CP_7983_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3166_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3166_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3166_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3166_sample_completed_
      -- 
    -- Element group sendModule_CP_7983_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3166_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3166_update_start_
      -- 
    -- Element group sendModule_CP_7983_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3166_update_completed__ps
      -- 
    sendModule_CP_7983_elements(32) <= sendModule_CP_7983_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3166_update_completed_
      -- 
    -- Element group sendModule_CP_7983_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => sendModule_CP_7983_elements(31), ack => sendModule_CP_7983_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_sample_start__ps
      -- CP-element group 34: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_Sample/req
      -- 
    req_8098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(34), ack => n_address1_3262_3167_buf_req_0); -- 
    -- Element group sendModule_CP_7983_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_update_start__ps
      -- CP-element group 35: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_update_start_
      -- CP-element group 35: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_Update/req
      -- 
    req_8103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(35), ack => n_address1_3262_3167_buf_req_1); -- 
    -- Element group sendModule_CP_7983_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_Sample/ack
      -- 
    ack_8099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_3262_3167_buf_ack_0, ack => sendModule_CP_7983_elements(36)); -- 
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address1_3167_Update/ack
      -- 
    ack_8104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_3262_3167_buf_ack_1, ack => sendModule_CP_7983_elements(37)); -- 
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	15 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	18 
    -- CP-element group 38: 	119 
    -- CP-element group 38: 	127 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	17 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_sample_start_
      -- 
    sendModule_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(18) & sendModule_CP_7983_elements(119) & sendModule_CP_7983_elements(127);
      gj_sendModule_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	15 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	138 
    -- CP-element group 39: 	292 
    -- CP-element group 39: 	300 
    -- CP-element group 39: 	308 
    -- CP-element group 39: 	316 
    -- CP-element group 39: 	340 
    -- CP-element group 39: 	348 
    -- CP-element group 39: 	324 
    -- CP-element group 39: 	332 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	19 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_update_start_
      -- 
    sendModule_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(138) & sendModule_CP_7983_elements(292) & sendModule_CP_7983_elements(300) & sendModule_CP_7983_elements(308) & sendModule_CP_7983_elements(316) & sendModule_CP_7983_elements(340) & sendModule_CP_7983_elements(348) & sendModule_CP_7983_elements(324) & sendModule_CP_7983_elements(332);
      gj_sendModule_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	17 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_sample_start__ps
      -- 
    sendModule_CP_7983_elements(40) <= sendModule_CP_7983_elements(17);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	18 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7983_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	19 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_update_start__ps
      -- 
    sendModule_CP_7983_elements(42) <= sendModule_CP_7983_elements(19);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	20 
    -- CP-element group 43: 	138 
    -- CP-element group 43: 	290 
    -- CP-element group 43: 	298 
    -- CP-element group 43: 	306 
    -- CP-element group 43: 	314 
    -- CP-element group 43: 	346 
    -- CP-element group 43: 	322 
    -- CP-element group 43: 	330 
    -- CP-element group 43: 	338 
    -- CP-element group 43:  members (15) 
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_update_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_resized_1
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_scaled_1
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_computed_1
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_resize_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_resize_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_resize_1/index_resize_req
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_resize_1/index_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_scale_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_scale_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_scale_1/scale_rename_req
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_index_scale_1/scale_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_final_index_sum_regn_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_final_index_sum_regn_Sample/req
      -- 
    req_8404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(43), ack => array_obj_ref_3294_index_offset_req_0); -- 
    -- Element group sendModule_CP_7983_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	13 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_loopback_trigger
      -- 
    sendModule_CP_7983_elements(44) <= sendModule_CP_7983_elements(13);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_loopback_sample_req
      -- CP-element group 45: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_loopback_sample_req_ps
      -- 
    phi_stmt_3168_loopback_sample_req_8115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3168_loopback_sample_req_8115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(45), ack => phi_stmt_3168_req_1); -- 
    -- Element group sendModule_CP_7983_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	14 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_entry_trigger
      -- 
    sendModule_CP_7983_elements(46) <= sendModule_CP_7983_elements(14);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_entry_sample_req
      -- CP-element group 47: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_entry_sample_req_ps
      -- 
    phi_stmt_3168_entry_sample_req_8118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3168_entry_sample_req_8118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(47), ack => phi_stmt_3168_req_0); -- 
    -- Element group sendModule_CP_7983_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_phi_mux_ack
      -- CP-element group 48: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3168_phi_mux_ack_ps
      -- 
    phi_stmt_3168_phi_mux_ack_8121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3168_ack_0, ack => sendModule_CP_7983_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_sample_start__ps
      -- 
    -- Element group sendModule_CP_7983_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_update_start__ps
      -- 
    -- Element group sendModule_CP_7983_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_Sample/rr
      -- 
    rr_8134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(51), ack => type_cast_3171_inst_req_0); -- 
    sendModule_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(49) & sendModule_CP_7983_elements(53);
      gj_sendModule_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_update_start_
      -- CP-element group 52: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_Update/cr
      -- 
    cr_8139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(52), ack => type_cast_3171_inst_req_1); -- 
    sendModule_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(50) & sendModule_CP_7983_elements(54);
      gj_sendModule_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_Sample/ra
      -- 
    ra_8135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3171_inst_ack_0, ack => sendModule_CP_7983_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3171_Update/ca
      -- 
    ca_8140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3171_inst_ack_1, ack => sendModule_CP_7983_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_sample_start__ps
      -- CP-element group 55: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_Sample/req
      -- 
    req_8152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(55), ack => n_address2_3276_3172_buf_req_0); -- 
    -- Element group sendModule_CP_7983_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_update_start__ps
      -- CP-element group 56: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_update_start_
      -- CP-element group 56: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_Update/req
      -- 
    req_8157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(56), ack => n_address2_3276_3172_buf_req_1); -- 
    -- Element group sendModule_CP_7983_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_sample_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_Sample/ack
      -- 
    ack_8153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_3276_3172_buf_ack_0, ack => sendModule_CP_7983_elements(57)); -- 
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_update_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_address2_3172_Update/ack
      -- 
    ack_8158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_3276_3172_buf_ack_1, ack => sendModule_CP_7983_elements(58)); -- 
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	15 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	18 
    -- CP-element group 59: 	119 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_sample_start_
      -- 
    sendModule_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(18) & sendModule_CP_7983_elements(119);
      gj_sendModule_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	15 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	64 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	19 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_update_start_
      -- 
    sendModule_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(64);
      gj_sendModule_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	17 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_sample_start__ps
      -- 
    sendModule_CP_7983_elements(61) <= sendModule_CP_7983_elements(17);
    -- CP-element group 62:  join  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	18 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7983_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	19 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_update_start__ps
      -- 
    sendModule_CP_7983_elements(63) <= sendModule_CP_7983_elements(19);
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	20 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	60 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_update_completed__ps
      -- 
    -- Element group sendModule_CP_7983_elements(64) is bound as output of CP function.
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	13 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_loopback_trigger
      -- 
    sendModule_CP_7983_elements(65) <= sendModule_CP_7983_elements(13);
    -- CP-element group 66:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_loopback_sample_req
      -- CP-element group 66: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_loopback_sample_req_ps
      -- 
    phi_stmt_3173_loopback_sample_req_8169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3173_loopback_sample_req_8169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(66), ack => phi_stmt_3173_req_1); -- 
    -- Element group sendModule_CP_7983_elements(66) is bound as output of CP function.
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	14 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_entry_trigger
      -- 
    sendModule_CP_7983_elements(67) <= sendModule_CP_7983_elements(14);
    -- CP-element group 68:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_entry_sample_req
      -- CP-element group 68: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_entry_sample_req_ps
      -- 
    phi_stmt_3173_entry_sample_req_8172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3173_entry_sample_req_8172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(68), ack => phi_stmt_3173_req_0); -- 
    -- Element group sendModule_CP_7983_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_phi_mux_ack
      -- CP-element group 69: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3173_phi_mux_ack_ps
      -- 
    phi_stmt_3173_phi_mux_ack_8175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3173_ack_0, ack => sendModule_CP_7983_elements(69)); -- 
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3176_sample_start__ps
      -- CP-element group 70: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3176_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3176_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3176_sample_completed_
      -- 
    -- Element group sendModule_CP_7983_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3176_update_start__ps
      -- CP-element group 71: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3176_update_start_
      -- 
    -- Element group sendModule_CP_7983_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3176_update_completed__ps
      -- 
    sendModule_CP_7983_elements(72) <= sendModule_CP_7983_elements(73);
    -- CP-element group 73:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	72 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3176_update_completed_
      -- 
    -- Element group sendModule_CP_7983_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => sendModule_CP_7983_elements(71), ack => sendModule_CP_7983_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_sample_start__ps
      -- CP-element group 74: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_Sample/req
      -- 
    req_8196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(74), ack => n_chl_3232_3177_buf_req_0); -- 
    -- Element group sendModule_CP_7983_elements(74) is bound as output of CP function.
    -- CP-element group 75:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_update_start__ps
      -- CP-element group 75: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_update_start_
      -- CP-element group 75: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_Update/req
      -- 
    req_8201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(75), ack => n_chl_3232_3177_buf_req_1); -- 
    -- Element group sendModule_CP_7983_elements(75) is bound as output of CP function.
    -- CP-element group 76:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_Sample/ack
      -- 
    ack_8197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3232_3177_buf_ack_0, ack => sendModule_CP_7983_elements(76)); -- 
    -- CP-element group 77:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_update_completed__ps
      -- CP-element group 77: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_chl_3177_Update/ack
      -- 
    ack_8202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3232_3177_buf_ack_1, ack => sendModule_CP_7983_elements(77)); -- 
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	15 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	18 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	17 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_sample_start_
      -- 
    sendModule_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(18);
      gj_sendModule_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	15 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	83 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	19 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_update_start_
      -- 
    sendModule_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(83);
      gj_sendModule_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_sample_start__ps
      -- 
    sendModule_CP_7983_elements(80) <= sendModule_CP_7983_elements(17);
    -- CP-element group 81:  join  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	18 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7983_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	19 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_update_start__ps
      -- 
    sendModule_CP_7983_elements(82) <= sendModule_CP_7983_elements(19);
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	20 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	79 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_update_completed__ps
      -- 
    -- Element group sendModule_CP_7983_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	13 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_loopback_trigger
      -- 
    sendModule_CP_7983_elements(84) <= sendModule_CP_7983_elements(13);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_loopback_sample_req
      -- CP-element group 85: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_loopback_sample_req_ps
      -- 
    phi_stmt_3178_loopback_sample_req_8213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3178_loopback_sample_req_8213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(85), ack => phi_stmt_3178_req_1); -- 
    -- Element group sendModule_CP_7983_elements(85) is bound as output of CP function.
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	14 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_entry_trigger
      -- 
    sendModule_CP_7983_elements(86) <= sendModule_CP_7983_elements(14);
    -- CP-element group 87:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_entry_sample_req
      -- CP-element group 87: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_entry_sample_req_ps
      -- 
    phi_stmt_3178_entry_sample_req_8216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3178_entry_sample_req_8216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(87), ack => phi_stmt_3178_req_0); -- 
    -- Element group sendModule_CP_7983_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_phi_mux_ack
      -- CP-element group 88: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3178_phi_mux_ack_ps
      -- 
    phi_stmt_3178_phi_mux_ack_8219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3178_ack_0, ack => sendModule_CP_7983_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3181_sample_start__ps
      -- CP-element group 89: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3181_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3181_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3181_sample_completed_
      -- 
    -- Element group sendModule_CP_7983_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3181_update_start__ps
      -- CP-element group 90: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3181_update_start_
      -- 
    -- Element group sendModule_CP_7983_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3181_update_completed__ps
      -- 
    sendModule_CP_7983_elements(91) <= sendModule_CP_7983_elements(92);
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	91 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3181_update_completed_
      -- 
    -- Element group sendModule_CP_7983_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => sendModule_CP_7983_elements(90), ack => sendModule_CP_7983_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_sample_start__ps
      -- CP-element group 93: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_Sample/req
      -- 
    req_8240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(93), ack => n_col_3213_3182_buf_req_0); -- 
    -- Element group sendModule_CP_7983_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_update_start__ps
      -- CP-element group 94: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_update_start_
      -- CP-element group 94: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_Update/req
      -- 
    req_8245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(94), ack => n_col_3213_3182_buf_req_1); -- 
    -- Element group sendModule_CP_7983_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_Sample/ack
      -- 
    ack_8241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3213_3182_buf_ack_0, ack => sendModule_CP_7983_elements(95)); -- 
    -- CP-element group 96:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_col_3182_Update/ack
      -- 
    ack_8246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3213_3182_buf_ack_1, ack => sendModule_CP_7983_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	15 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	18 
    -- CP-element group 97: 	119 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	17 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_sample_start_
      -- 
    sendModule_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(18) & sendModule_CP_7983_elements(119);
      gj_sendModule_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	15 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	102 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	19 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_update_start_
      -- 
    sendModule_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(102);
      gj_sendModule_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	17 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_sample_start__ps
      -- 
    sendModule_CP_7983_elements(99) <= sendModule_CP_7983_elements(17);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	18 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7983_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	19 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_update_start__ps
      -- 
    sendModule_CP_7983_elements(101) <= sendModule_CP_7983_elements(19);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	20 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	98 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_update_completed__ps
      -- 
    -- Element group sendModule_CP_7983_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	13 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_loopback_trigger
      -- 
    sendModule_CP_7983_elements(103) <= sendModule_CP_7983_elements(13);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_loopback_sample_req
      -- CP-element group 104: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_loopback_sample_req_ps
      -- 
    phi_stmt_3183_loopback_sample_req_8257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3183_loopback_sample_req_8257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(104), ack => phi_stmt_3183_req_1); -- 
    -- Element group sendModule_CP_7983_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	14 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_entry_trigger
      -- 
    sendModule_CP_7983_elements(105) <= sendModule_CP_7983_elements(14);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_entry_sample_req
      -- CP-element group 106: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_entry_sample_req_ps
      -- 
    phi_stmt_3183_entry_sample_req_8260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3183_entry_sample_req_8260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(106), ack => phi_stmt_3183_req_0); -- 
    -- Element group sendModule_CP_7983_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_phi_mux_ack
      -- CP-element group 107: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/phi_stmt_3183_phi_mux_ack_ps
      -- 
    phi_stmt_3183_phi_mux_ack_8263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3183_ack_0, ack => sendModule_CP_7983_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3186_sample_start__ps
      -- CP-element group 108: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3186_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3186_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3186_sample_completed_
      -- 
    -- Element group sendModule_CP_7983_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3186_update_start__ps
      -- CP-element group 109: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3186_update_start_
      -- 
    -- Element group sendModule_CP_7983_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3186_update_completed__ps
      -- 
    sendModule_CP_7983_elements(110) <= sendModule_CP_7983_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3186_update_completed_
      -- 
    -- Element group sendModule_CP_7983_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => sendModule_CP_7983_elements(109), ack => sendModule_CP_7983_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_sample_start__ps
      -- CP-element group 112: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_Sample/req
      -- 
    req_8284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(112), ack => n_row_3224_3187_buf_req_0); -- 
    -- Element group sendModule_CP_7983_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_update_start__ps
      -- CP-element group 113: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_update_start_
      -- CP-element group 113: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_Update/req
      -- 
    req_8289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(113), ack => n_row_3224_3187_buf_req_1); -- 
    -- Element group sendModule_CP_7983_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_Sample/ack
      -- 
    ack_8285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3224_3187_buf_ack_0, ack => sendModule_CP_7983_elements(114)); -- 
    -- CP-element group 115:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_update_completed__ps
      -- CP-element group 115: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/R_n_row_3187_Update/ack
      -- 
    ack_8290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3224_3187_buf_ack_1, ack => sendModule_CP_7983_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	15 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_Sample/rr
      -- 
    rr_8299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(116), ack => SUB_u16_u16_3197_inst_req_0); -- 
    sendModule_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(118);
      gj_sendModule_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	18 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_update_start_
      -- CP-element group 117: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_Update/cr
      -- 
    cr_8304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(117), ack => SUB_u16_u16_3197_inst_req_1); -- 
    sendModule_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(18) & sendModule_CP_7983_elements(119);
      gj_sendModule_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_Sample/ra
      -- 
    ra_8300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3197_inst_ack_0, ack => sendModule_CP_7983_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	16 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	21 
    -- CP-element group 119: 	38 
    -- CP-element group 119: 	59 
    -- CP-element group 119: 	97 
    -- CP-element group 119: 	117 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3197_Update/ca
      -- 
    ca_8305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3197_inst_ack_1, ack => sendModule_CP_7983_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	15 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_Sample/rr
      -- 
    rr_8313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(120), ack => type_cast_3235_inst_req_0); -- 
    sendModule_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(122);
      gj_sendModule_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	18 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_update_start_
      -- CP-element group 121: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_Update/cr
      -- 
    cr_8318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(121), ack => type_cast_3235_inst_req_1); -- 
    sendModule_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(18) & sendModule_CP_7983_elements(123);
      gj_sendModule_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_Sample/ra
      -- 
    ra_8314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3235_inst_ack_0, ack => sendModule_CP_7983_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	386 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	21 
    -- CP-element group 123: 	121 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3235_Update/ca
      -- 
    ca_8319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3235_inst_ack_1, ack => sendModule_CP_7983_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	15 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_Sample/rr
      -- 
    rr_8327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(124), ack => type_cast_3244_inst_req_0); -- 
    sendModule_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(126);
      gj_sendModule_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	18 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_update_start_
      -- CP-element group 125: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_Update/$entry
      -- CP-element group 125: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_Update/cr
      -- 
    cr_8332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(125), ack => type_cast_3244_inst_req_1); -- 
    sendModule_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(18) & sendModule_CP_7983_elements(127);
      gj_sendModule_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_Sample/ra
      -- 
    ra_8328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3244_inst_ack_0, ack => sendModule_CP_7983_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	386 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	38 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/type_cast_3244_Update/ca
      -- 
    ca_8333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3244_inst_ack_1, ack => sendModule_CP_7983_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	132 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	133 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	133 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_request/$entry
      -- CP-element group 128: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_request/req
      -- 
    req_8373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(128), ack => addr_of_3285_final_reg_req_0); -- 
    sendModule_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(132) & sendModule_CP_7983_elements(133);
      gj_sendModule_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	15 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	144 
    -- CP-element group 129: 	356 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	134 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_update_start_
      -- CP-element group 129: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_complete/$entry
      -- CP-element group 129: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_complete/req
      -- 
    req_8378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(129), ack => addr_of_3285_final_reg_req_1); -- 
    sendModule_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(144) & sendModule_CP_7983_elements(356);
      gj_sendModule_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	15 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	133 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_final_index_sum_regn_update_start
      -- CP-element group 130: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_final_index_sum_regn_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_final_index_sum_regn_Update/req
      -- 
    req_8363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(130), ack => array_obj_ref_3284_index_offset_req_1); -- 
    sendModule_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(133);
      gj_sendModule_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	24 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	386 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	22 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_final_index_sum_regn_sample_complete
      -- CP-element group 131: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_final_index_sum_regn_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_final_index_sum_regn_Sample/ack
      -- 
    ack_8359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3284_index_offset_ack_0, ack => sendModule_CP_7983_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	128 
    -- CP-element group 132:  members (8) 
      -- CP-element group 132: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_root_address_calculated
      -- CP-element group 132: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_offset_calculated
      -- CP-element group 132: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_final_index_sum_regn_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_final_index_sum_regn_Update/ack
      -- CP-element group 132: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_base_plus_offset/$entry
      -- CP-element group 132: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_base_plus_offset/$exit
      -- CP-element group 132: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_base_plus_offset/sum_rename_req
      -- CP-element group 132: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3284_base_plus_offset/sum_rename_ack
      -- 
    ack_8364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3284_index_offset_ack_1, ack => sendModule_CP_7983_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	128 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	128 
    -- CP-element group 133: 	130 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_request/$exit
      -- CP-element group 133: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_request/ack
      -- 
    ack_8374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3285_final_reg_ack_0, ack => sendModule_CP_7983_elements(133)); -- 
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	129 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	142 
    -- CP-element group 134: 	354 
    -- CP-element group 134:  members (19) 
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_complete/$exit
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3285_complete/ack
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_base_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_word_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_root_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_base_address_resized
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_base_addr_resize/$entry
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_base_addr_resize/$exit
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_base_addr_resize/base_resize_req
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_base_addr_resize/base_resize_ack
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_base_plus_offset/$entry
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_base_plus_offset/$exit
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_base_plus_offset/sum_rename_req
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_base_plus_offset/sum_rename_ack
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_word_addrgen/$entry
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_word_addrgen/$exit
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_word_addrgen/root_register_req
      -- CP-element group 134: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_word_addrgen/root_register_ack
      -- 
    ack_8379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3285_final_reg_ack_1, ack => sendModule_CP_7983_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	139 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	140 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	140 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_request/$entry
      -- CP-element group 135: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_request/req
      -- 
    req_8419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(135), ack => addr_of_3295_final_reg_req_0); -- 
    sendModule_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(139) & sendModule_CP_7983_elements(140);
      gj_sendModule_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	15 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	368 
    -- CP-element group 136: 	148 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	141 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_update_start_
      -- CP-element group 136: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_complete/req
      -- 
    req_8424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(136), ack => addr_of_3295_final_reg_req_1); -- 
    sendModule_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(368) & sendModule_CP_7983_elements(148);
      gj_sendModule_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	15 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	140 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_final_index_sum_regn_update_start
      -- CP-element group 137: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_final_index_sum_regn_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_final_index_sum_regn_Update/req
      -- 
    req_8409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(137), ack => array_obj_ref_3294_index_offset_req_1); -- 
    sendModule_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(140);
      gj_sendModule_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	43 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	386 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	39 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_final_index_sum_regn_sample_complete
      -- CP-element group 138: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_final_index_sum_regn_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_final_index_sum_regn_Sample/ack
      -- 
    ack_8405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3294_index_offset_ack_0, ack => sendModule_CP_7983_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	135 
    -- CP-element group 139:  members (8) 
      -- CP-element group 139: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_offset_calculated
      -- CP-element group 139: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_final_index_sum_regn_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_final_index_sum_regn_Update/ack
      -- CP-element group 139: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_base_plus_offset/$entry
      -- CP-element group 139: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_base_plus_offset/$exit
      -- CP-element group 139: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_base_plus_offset/sum_rename_req
      -- CP-element group 139: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/array_obj_ref_3294_base_plus_offset/sum_rename_ack
      -- 
    ack_8410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3294_index_offset_ack_1, ack => sendModule_CP_7983_elements(139)); -- 
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	135 
    -- CP-element group 140: successors 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	137 
    -- CP-element group 140: 	135 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_request/$exit
      -- CP-element group 140: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_request/ack
      -- 
    ack_8420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3295_final_reg_ack_0, ack => sendModule_CP_7983_elements(140)); -- 
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	136 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	146 
    -- CP-element group 141: 	366 
    -- CP-element group 141:  members (19) 
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_base_address_resized
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_word_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_word_addrgen/$exit
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_word_addrgen/root_register_ack
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_word_addrgen/root_register_req
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_base_addr_resize/base_resize_ack
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_base_addr_resize/base_resize_req
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_base_addr_resize/$exit
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_base_addr_resize/$entry
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_word_addrgen/$entry
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_complete/$exit
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/addr_of_3295_complete/ack
      -- CP-element group 141: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_base_address_calculated
      -- 
    ack_8425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3295_final_reg_ack_1, ack => sendModule_CP_7983_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	134 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	376 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (5) 
      -- CP-element group 142: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Sample/word_access_start/$entry
      -- CP-element group 142: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Sample/word_access_start/word_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Sample/word_access_start/word_0/rr
      -- 
    rr_8458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(142), ack => ptr_deref_3299_load_0_req_0); -- 
    sendModule_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(134) & sendModule_CP_7983_elements(376);
      gj_sendModule_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	164 
    -- CP-element group 143: 	168 
    -- CP-element group 143: 	172 
    -- CP-element group 143: 	176 
    -- CP-element group 143: 	180 
    -- CP-element group 143: 	184 
    -- CP-element group 143: 	188 
    -- CP-element group 143: 	192 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_update_start_
      -- CP-element group 143: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/word_access_complete/$entry
      -- CP-element group 143: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/word_access_complete/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/word_access_complete/word_0/cr
      -- 
    cr_8469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(143), ack => ptr_deref_3299_load_0_req_1); -- 
    sendModule_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(164) & sendModule_CP_7983_elements(168) & sendModule_CP_7983_elements(172) & sendModule_CP_7983_elements(176) & sendModule_CP_7983_elements(180) & sendModule_CP_7983_elements(184) & sendModule_CP_7983_elements(188) & sendModule_CP_7983_elements(192);
      gj_sendModule_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	383 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	129 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Sample/word_access_start/word_0/ra
      -- 
    ra_8459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3299_load_0_ack_0, ack => sendModule_CP_7983_elements(144)); -- 
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	166 
    -- CP-element group 145: 	170 
    -- CP-element group 145: 	174 
    -- CP-element group 145: 	178 
    -- CP-element group 145: 	182 
    -- CP-element group 145: 	186 
    -- CP-element group 145: 	190 
    -- CP-element group 145: 	162 
    -- CP-element group 145:  members (9) 
      -- CP-element group 145: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/word_access_complete/word_0/ca
      -- CP-element group 145: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/ptr_deref_3299_Merge/$entry
      -- CP-element group 145: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/ptr_deref_3299_Merge/$exit
      -- CP-element group 145: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/ptr_deref_3299_Merge/merge_req
      -- CP-element group 145: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_Update/ptr_deref_3299_Merge/merge_ack
      -- 
    ca_8470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3299_load_0_ack_1, ack => sendModule_CP_7983_elements(145)); -- 
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	141 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	376 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Sample/word_access_start/word_0/$entry
      -- CP-element group 146: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Sample/word_access_start/word_0/rr
      -- CP-element group 146: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Sample/word_access_start/$entry
      -- CP-element group 146: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_sample_start_
      -- 
    rr_8508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(146), ack => ptr_deref_3303_load_0_req_0); -- 
    sendModule_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(141) & sendModule_CP_7983_elements(376);
      gj_sendModule_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	196 
    -- CP-element group 147: 	200 
    -- CP-element group 147: 	204 
    -- CP-element group 147: 	208 
    -- CP-element group 147: 	212 
    -- CP-element group 147: 	216 
    -- CP-element group 147: 	220 
    -- CP-element group 147: 	224 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/word_access_complete/$entry
      -- CP-element group 147: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/word_access_complete/word_0/cr
      -- CP-element group 147: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/word_access_complete/word_0/$entry
      -- CP-element group 147: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_update_start_
      -- 
    cr_8519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(147), ack => ptr_deref_3303_load_0_req_1); -- 
    sendModule_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(196) & sendModule_CP_7983_elements(200) & sendModule_CP_7983_elements(204) & sendModule_CP_7983_elements(208) & sendModule_CP_7983_elements(212) & sendModule_CP_7983_elements(216) & sendModule_CP_7983_elements(220) & sendModule_CP_7983_elements(224);
      gj_sendModule_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	384 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	136 
    -- CP-element group 148:  members (5) 
      -- CP-element group 148: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Sample/word_access_start/word_0/ra
      -- CP-element group 148: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Sample/word_access_start/word_0/$exit
      -- CP-element group 148: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Sample/word_access_start/$exit
      -- CP-element group 148: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_sample_completed_
      -- 
    ra_8509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3303_load_0_ack_0, ack => sendModule_CP_7983_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	194 
    -- CP-element group 149: 	198 
    -- CP-element group 149: 	202 
    -- CP-element group 149: 	206 
    -- CP-element group 149: 	210 
    -- CP-element group 149: 	214 
    -- CP-element group 149: 	218 
    -- CP-element group 149: 	222 
    -- CP-element group 149:  members (9) 
      -- CP-element group 149: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/word_access_complete/$exit
      -- CP-element group 149: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/word_access_complete/word_0/$exit
      -- CP-element group 149: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/ptr_deref_3303_Merge/$exit
      -- CP-element group 149: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/ptr_deref_3303_Merge/merge_ack
      -- CP-element group 149: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/ptr_deref_3303_Merge/merge_req
      -- CP-element group 149: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/ptr_deref_3303_Merge/$entry
      -- CP-element group 149: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_Update/word_access_complete/word_0/ca
      -- CP-element group 149: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_update_completed_
      -- 
    ca_8520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3303_load_0_ack_1, ack => sendModule_CP_7983_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	15 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_sample_start_
      -- 
    rr_8533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(150), ack => RPIPE_output_pipe_3306_inst_req_0); -- 
    sendModule_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(153);
      gj_sendModule_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	156 
    -- CP-element group 151: 	160 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_update_start_
      -- CP-element group 151: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_Update/cr
      -- 
    cr_8538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(151), ack => RPIPE_output_pipe_3306_inst_req_1); -- 
    sendModule_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(152) & sendModule_CP_7983_elements(156) & sendModule_CP_7983_elements(160);
      gj_sendModule_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	151 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_sample_completed_
      -- 
    ra_8534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3306_inst_ack_0, ack => sendModule_CP_7983_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	158 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/RPIPE_output_pipe_3306_Update/ca
      -- 
    ca_8539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3306_inst_ack_1, ack => sendModule_CP_7983_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_Sample/$entry
      -- 
    rr_8547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(154), ack => slice_3310_inst_req_0); -- 
    sendModule_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(153) & sendModule_CP_7983_elements(156);
      gj_sendModule_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	272 
    -- CP-element group 155: 	280 
    -- CP-element group 155: 	288 
    -- CP-element group 155: 	256 
    -- CP-element group 155: 	264 
    -- CP-element group 155: 	232 
    -- CP-element group 155: 	240 
    -- CP-element group 155: 	248 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_update_start_
      -- CP-element group 155: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_Update/cr
      -- 
    cr_8552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(155), ack => slice_3310_inst_req_1); -- 
    sendModule_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(272) & sendModule_CP_7983_elements(280) & sendModule_CP_7983_elements(288) & sendModule_CP_7983_elements(256) & sendModule_CP_7983_elements(264) & sendModule_CP_7983_elements(232) & sendModule_CP_7983_elements(240) & sendModule_CP_7983_elements(248);
      gj_sendModule_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	151 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_sample_completed_
      -- 
    ra_8548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3310_inst_ack_0, ack => sendModule_CP_7983_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	270 
    -- CP-element group 157: 	278 
    -- CP-element group 157: 	286 
    -- CP-element group 157: 	254 
    -- CP-element group 157: 	262 
    -- CP-element group 157: 	238 
    -- CP-element group 157: 	246 
    -- CP-element group 157: 	230 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3310_Update/ca
      -- 
    ca_8553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3310_inst_ack_1, ack => sendModule_CP_7983_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	153 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_Sample/rr
      -- 
    rr_8561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(158), ack => slice_3314_inst_req_0); -- 
    sendModule_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(153) & sendModule_CP_7983_elements(160);
      gj_sendModule_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	296 
    -- CP-element group 159: 	304 
    -- CP-element group 159: 	312 
    -- CP-element group 159: 	320 
    -- CP-element group 159: 	344 
    -- CP-element group 159: 	352 
    -- CP-element group 159: 	328 
    -- CP-element group 159: 	336 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_update_start_
      -- CP-element group 159: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_Update/cr
      -- CP-element group 159: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_Update/$entry
      -- 
    cr_8566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(159), ack => slice_3314_inst_req_1); -- 
    sendModule_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(296) & sendModule_CP_7983_elements(304) & sendModule_CP_7983_elements(312) & sendModule_CP_7983_elements(320) & sendModule_CP_7983_elements(344) & sendModule_CP_7983_elements(352) & sendModule_CP_7983_elements(328) & sendModule_CP_7983_elements(336);
      gj_sendModule_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	151 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_Sample/ra
      -- 
    ra_8562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3314_inst_ack_0, ack => sendModule_CP_7983_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	294 
    -- CP-element group 161: 	302 
    -- CP-element group 161: 	310 
    -- CP-element group 161: 	318 
    -- CP-element group 161: 	342 
    -- CP-element group 161: 	350 
    -- CP-element group 161: 	326 
    -- CP-element group 161: 	334 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_Update/ca
      -- CP-element group 161: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3314_Update/$exit
      -- 
    ca_8567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3314_inst_ack_1, ack => sendModule_CP_7983_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	145 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_Sample/rr
      -- 
    rr_8575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(162), ack => slice_3318_inst_req_0); -- 
    sendModule_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(145) & sendModule_CP_7983_elements(164);
      gj_sendModule_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	360 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_Update/cr
      -- 
    cr_8580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(163), ack => slice_3318_inst_req_1); -- 
    sendModule_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	143 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_Sample/ra
      -- 
    ra_8576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3318_inst_ack_0, ack => sendModule_CP_7983_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	358 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3318_Update/ca
      -- 
    ca_8581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3318_inst_ack_1, ack => sendModule_CP_7983_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	145 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_Sample/rr
      -- 
    rr_8589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(166), ack => slice_3322_inst_req_0); -- 
    sendModule_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(145) & sendModule_CP_7983_elements(168);
      gj_sendModule_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	360 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_update_start_
      -- CP-element group 167: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_Update/cr
      -- 
    cr_8594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(167), ack => slice_3322_inst_req_1); -- 
    sendModule_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: 	143 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_Sample/ra
      -- 
    ra_8590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3322_inst_ack_0, ack => sendModule_CP_7983_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	358 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3322_Update/ca
      -- 
    ca_8595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3322_inst_ack_1, ack => sendModule_CP_7983_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	145 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_Sample/rr
      -- 
    rr_8603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(170), ack => slice_3326_inst_req_0); -- 
    sendModule_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(145) & sendModule_CP_7983_elements(172);
      gj_sendModule_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	360 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_update_start_
      -- CP-element group 171: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_Update/cr
      -- 
    cr_8608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(171), ack => slice_3326_inst_req_1); -- 
    sendModule_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: 	143 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_Sample/ra
      -- 
    ra_8604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3326_inst_ack_0, ack => sendModule_CP_7983_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	358 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3326_Update/ca
      -- 
    ca_8609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3326_inst_ack_1, ack => sendModule_CP_7983_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	145 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_Sample/rr
      -- 
    rr_8617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(174), ack => slice_3330_inst_req_0); -- 
    sendModule_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(145) & sendModule_CP_7983_elements(176);
      gj_sendModule_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	360 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_update_start_
      -- CP-element group 175: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_Update/cr
      -- 
    cr_8622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(175), ack => slice_3330_inst_req_1); -- 
    sendModule_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: 	143 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_Sample/ra
      -- 
    ra_8618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3330_inst_ack_0, ack => sendModule_CP_7983_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	358 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3330_Update/ca
      -- 
    ca_8623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3330_inst_ack_1, ack => sendModule_CP_7983_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	145 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_Sample/rr
      -- 
    rr_8631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(178), ack => slice_3334_inst_req_0); -- 
    sendModule_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(145) & sendModule_CP_7983_elements(180);
      gj_sendModule_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	360 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_update_start_
      -- CP-element group 179: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_Update/cr
      -- 
    cr_8636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(179), ack => slice_3334_inst_req_1); -- 
    sendModule_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	143 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_Sample/ra
      -- 
    ra_8632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3334_inst_ack_0, ack => sendModule_CP_7983_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	358 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3334_Update/ca
      -- 
    ca_8637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3334_inst_ack_1, ack => sendModule_CP_7983_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	145 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_Sample/rr
      -- 
    rr_8645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(182), ack => slice_3338_inst_req_0); -- 
    sendModule_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(145) & sendModule_CP_7983_elements(184);
      gj_sendModule_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	360 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_update_start_
      -- CP-element group 183: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_Update/cr
      -- 
    cr_8650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(183), ack => slice_3338_inst_req_1); -- 
    sendModule_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	143 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_Sample/ra
      -- 
    ra_8646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3338_inst_ack_0, ack => sendModule_CP_7983_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	358 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3338_Update/ca
      -- 
    ca_8651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3338_inst_ack_1, ack => sendModule_CP_7983_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	145 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_Sample/rr
      -- 
    rr_8659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(186), ack => slice_3342_inst_req_0); -- 
    sendModule_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(145) & sendModule_CP_7983_elements(188);
      gj_sendModule_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	360 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_update_start_
      -- CP-element group 187: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_Update/cr
      -- 
    cr_8664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(187), ack => slice_3342_inst_req_1); -- 
    sendModule_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	143 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_Sample/ra
      -- 
    ra_8660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3342_inst_ack_0, ack => sendModule_CP_7983_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	358 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3342_Update/ca
      -- 
    ca_8665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3342_inst_ack_1, ack => sendModule_CP_7983_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	145 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_Sample/rr
      -- 
    rr_8673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(190), ack => slice_3346_inst_req_0); -- 
    sendModule_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(145) & sendModule_CP_7983_elements(192);
      gj_sendModule_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	360 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_update_start_
      -- CP-element group 191: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_Update/cr
      -- 
    cr_8678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(191), ack => slice_3346_inst_req_1); -- 
    sendModule_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	143 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_Sample/ra
      -- 
    ra_8674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3346_inst_ack_0, ack => sendModule_CP_7983_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	358 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3346_Update/ca
      -- 
    ca_8679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3346_inst_ack_1, ack => sendModule_CP_7983_elements(193)); -- 
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	149 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_Sample/rr
      -- 
    rr_8687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(194), ack => slice_3350_inst_req_0); -- 
    sendModule_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(149) & sendModule_CP_7983_elements(196);
      gj_sendModule_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	372 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_update_start_
      -- CP-element group 195: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_Update/cr
      -- 
    cr_8692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(195), ack => slice_3350_inst_req_1); -- 
    sendModule_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	147 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_Sample/ra
      -- 
    ra_8688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3350_inst_ack_0, ack => sendModule_CP_7983_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	370 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3350_Update/ca
      -- 
    ca_8693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3350_inst_ack_1, ack => sendModule_CP_7983_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	149 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_Sample/rr
      -- 
    rr_8701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(198), ack => slice_3354_inst_req_0); -- 
    sendModule_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(149) & sendModule_CP_7983_elements(200);
      gj_sendModule_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	372 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_update_start_
      -- CP-element group 199: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_Update/cr
      -- 
    cr_8706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(199), ack => slice_3354_inst_req_1); -- 
    sendModule_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	147 
    -- CP-element group 200: 	198 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_Sample/ra
      -- 
    ra_8702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3354_inst_ack_0, ack => sendModule_CP_7983_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	370 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3354_Update/ca
      -- 
    ca_8707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3354_inst_ack_1, ack => sendModule_CP_7983_elements(201)); -- 
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	149 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_Sample/rr
      -- 
    rr_8715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(202), ack => slice_3358_inst_req_0); -- 
    sendModule_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(149) & sendModule_CP_7983_elements(204);
      gj_sendModule_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	372 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_update_start_
      -- CP-element group 203: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_Update/cr
      -- 
    cr_8720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(203), ack => slice_3358_inst_req_1); -- 
    sendModule_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	147 
    -- CP-element group 204: 	202 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_Sample/ra
      -- 
    ra_8716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3358_inst_ack_0, ack => sendModule_CP_7983_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	370 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3358_Update/ca
      -- 
    ca_8721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3358_inst_ack_1, ack => sendModule_CP_7983_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	149 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_Sample/rr
      -- 
    rr_8729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(206), ack => slice_3362_inst_req_0); -- 
    sendModule_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(149) & sendModule_CP_7983_elements(208);
      gj_sendModule_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	372 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_update_start_
      -- CP-element group 207: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_Update/cr
      -- 
    cr_8734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(207), ack => slice_3362_inst_req_1); -- 
    sendModule_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	147 
    -- CP-element group 208: 	206 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_Sample/ra
      -- 
    ra_8730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3362_inst_ack_0, ack => sendModule_CP_7983_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	370 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3362_Update/ca
      -- 
    ca_8735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3362_inst_ack_1, ack => sendModule_CP_7983_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	149 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_Sample/rr
      -- 
    rr_8743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(210), ack => slice_3366_inst_req_0); -- 
    sendModule_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(149) & sendModule_CP_7983_elements(212);
      gj_sendModule_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	372 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_update_start_
      -- CP-element group 211: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_Update/cr
      -- 
    cr_8748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(211), ack => slice_3366_inst_req_1); -- 
    sendModule_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	147 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_Sample/ra
      -- 
    ra_8744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3366_inst_ack_0, ack => sendModule_CP_7983_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	370 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3366_Update/ca
      -- 
    ca_8749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3366_inst_ack_1, ack => sendModule_CP_7983_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	149 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_Sample/rr
      -- 
    rr_8757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(214), ack => slice_3370_inst_req_0); -- 
    sendModule_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(149) & sendModule_CP_7983_elements(216);
      gj_sendModule_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	372 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_update_start_
      -- CP-element group 215: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_Update/cr
      -- 
    cr_8762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(215), ack => slice_3370_inst_req_1); -- 
    sendModule_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	147 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_Sample/ra
      -- 
    ra_8758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3370_inst_ack_0, ack => sendModule_CP_7983_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	370 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3370_Update/ca
      -- 
    ca_8763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3370_inst_ack_1, ack => sendModule_CP_7983_elements(217)); -- 
    -- CP-element group 218:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	149 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_Sample/rr
      -- 
    rr_8771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(218), ack => slice_3374_inst_req_0); -- 
    sendModule_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(149) & sendModule_CP_7983_elements(220);
      gj_sendModule_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: marked-predecessors 
    -- CP-element group 219: 	372 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_update_start_
      -- CP-element group 219: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_Update/cr
      -- 
    cr_8776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(219), ack => slice_3374_inst_req_1); -- 
    sendModule_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	147 
    -- CP-element group 220: 	218 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_Sample/ra
      -- 
    ra_8772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3374_inst_ack_0, ack => sendModule_CP_7983_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	370 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3374_Update/ca
      -- 
    ca_8777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3374_inst_ack_1, ack => sendModule_CP_7983_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	149 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_Sample/rr
      -- 
    rr_8785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(222), ack => slice_3378_inst_req_0); -- 
    sendModule_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(149) & sendModule_CP_7983_elements(224);
      gj_sendModule_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	372 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_update_start_
      -- CP-element group 223: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_Update/cr
      -- 
    cr_8790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(223), ack => slice_3378_inst_req_1); -- 
    sendModule_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	147 
    -- CP-element group 224: 	222 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_Sample/ra
      -- 
    ra_8786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3378_inst_ack_0, ack => sendModule_CP_7983_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	370 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/slice_3378_Update/ca
      -- 
    ca_8791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3378_inst_ack_1, ack => sendModule_CP_7983_elements(225)); -- 
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	24 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_Sample/rr
      -- 
    rr_8799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(226), ack => EQ_u3_u1_3391_inst_req_0); -- 
    sendModule_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(24) & sendModule_CP_7983_elements(228);
      gj_sendModule_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	360 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_update_start_
      -- CP-element group 227: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_Update/cr
      -- 
    cr_8804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(227), ack => EQ_u3_u1_3391_inst_req_1); -- 
    sendModule_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	22 
    -- CP-element group 228: 	226 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_Sample/ra
      -- 
    ra_8800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3391_inst_ack_0, ack => sendModule_CP_7983_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	358 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3391_Update/ca
      -- 
    ca_8805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3391_inst_ack_1, ack => sendModule_CP_7983_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	157 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_Sample/req
      -- 
    req_8813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(230), ack => W_output_data1_3266_delayed_13_0_3393_inst_req_0); -- 
    sendModule_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(157) & sendModule_CP_7983_elements(232);
      gj_sendModule_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: marked-predecessors 
    -- CP-element group 231: 	360 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	233 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_update_start_
      -- CP-element group 231: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_Update/req
      -- 
    req_8818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(231), ack => W_output_data1_3266_delayed_13_0_3393_inst_req_1); -- 
    sendModule_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: 	155 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_Sample/ack
      -- 
    ack_8814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3266_delayed_13_0_3393_inst_ack_0, ack => sendModule_CP_7983_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	231 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	358 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3395_Update/ack
      -- 
    ack_8819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3266_delayed_13_0_3393_inst_ack_1, ack => sendModule_CP_7983_elements(233)); -- 
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	24 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_Sample/rr
      -- 
    rr_8827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(234), ack => EQ_u3_u1_3405_inst_req_0); -- 
    sendModule_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(24) & sendModule_CP_7983_elements(236);
      gj_sendModule_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: marked-predecessors 
    -- CP-element group 235: 	360 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_update_start_
      -- CP-element group 235: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_Update/cr
      -- 
    cr_8832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(235), ack => EQ_u3_u1_3405_inst_req_1); -- 
    sendModule_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	22 
    -- CP-element group 236: 	234 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_Sample/ra
      -- 
    ra_8828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3405_inst_ack_0, ack => sendModule_CP_7983_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	358 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3405_Update/ca
      -- 
    ca_8833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3405_inst_ack_1, ack => sendModule_CP_7983_elements(237)); -- 
    -- CP-element group 238:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	157 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_Sample/req
      -- 
    req_8841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(238), ack => W_output_data1_3274_delayed_13_0_3407_inst_req_0); -- 
    sendModule_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(157) & sendModule_CP_7983_elements(240);
      gj_sendModule_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: marked-predecessors 
    -- CP-element group 239: 	360 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_update_start_
      -- CP-element group 239: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_Update/req
      -- 
    req_8846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(239), ack => W_output_data1_3274_delayed_13_0_3407_inst_req_1); -- 
    sendModule_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: 	155 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_sample_completed_
      -- CP-element group 240: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_Sample/ack
      -- 
    ack_8842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3274_delayed_13_0_3407_inst_ack_0, ack => sendModule_CP_7983_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	358 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_update_completed_
      -- CP-element group 241: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3409_Update/ack
      -- 
    ack_8847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3274_delayed_13_0_3407_inst_ack_1, ack => sendModule_CP_7983_elements(241)); -- 
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	24 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	244 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_Sample/rr
      -- 
    rr_8855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(242), ack => EQ_u3_u1_3419_inst_req_0); -- 
    sendModule_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(24) & sendModule_CP_7983_elements(244);
      gj_sendModule_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: marked-predecessors 
    -- CP-element group 243: 	360 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	245 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_update_start_
      -- CP-element group 243: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_Update/cr
      -- 
    cr_8860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(243), ack => EQ_u3_u1_3419_inst_req_1); -- 
    sendModule_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_243 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	22 
    -- CP-element group 244: 	242 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_Sample/ra
      -- 
    ra_8856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3419_inst_ack_0, ack => sendModule_CP_7983_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	243 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	358 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3419_Update/ca
      -- 
    ca_8861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3419_inst_ack_1, ack => sendModule_CP_7983_elements(245)); -- 
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	157 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	248 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_Sample/req
      -- 
    req_8869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(246), ack => W_output_data1_3282_delayed_13_0_3421_inst_req_0); -- 
    sendModule_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(157) & sendModule_CP_7983_elements(248);
      gj_sendModule_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: marked-predecessors 
    -- CP-element group 247: 	360 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	249 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_update_start_
      -- CP-element group 247: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_Update/req
      -- 
    req_8874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(247), ack => W_output_data1_3282_delayed_13_0_3421_inst_req_1); -- 
    sendModule_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: 	155 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_Sample/ack
      -- 
    ack_8870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3282_delayed_13_0_3421_inst_ack_0, ack => sendModule_CP_7983_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	358 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3423_Update/ack
      -- 
    ack_8875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3282_delayed_13_0_3421_inst_ack_1, ack => sendModule_CP_7983_elements(249)); -- 
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	24 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	252 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_Sample/rr
      -- 
    rr_8883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(250), ack => EQ_u3_u1_3433_inst_req_0); -- 
    sendModule_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(24) & sendModule_CP_7983_elements(252);
      gj_sendModule_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: marked-predecessors 
    -- CP-element group 251: 	360 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	253 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_update_start_
      -- CP-element group 251: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_Update/cr
      -- 
    cr_8888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(251), ack => EQ_u3_u1_3433_inst_req_1); -- 
    sendModule_cp_element_group_251: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_251"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_251 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(251), clk => clk, reset => reset); --
    end block;
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	22 
    -- CP-element group 252: 	250 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_Sample/ra
      -- 
    ra_8884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3433_inst_ack_0, ack => sendModule_CP_7983_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	251 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	358 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3433_Update/ca
      -- 
    ca_8889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3433_inst_ack_1, ack => sendModule_CP_7983_elements(253)); -- 
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	157 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_Sample/req
      -- 
    req_8897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(254), ack => W_output_data1_3290_delayed_13_0_3435_inst_req_0); -- 
    sendModule_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(157) & sendModule_CP_7983_elements(256);
      gj_sendModule_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: marked-predecessors 
    -- CP-element group 255: 	360 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_update_start_
      -- CP-element group 255: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_Update/req
      -- 
    req_8902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(255), ack => W_output_data1_3290_delayed_13_0_3435_inst_req_1); -- 
    sendModule_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: marked-successors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: 	155 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_Sample/ack
      -- 
    ack_8898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3290_delayed_13_0_3435_inst_ack_0, ack => sendModule_CP_7983_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	358 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3437_Update/ack
      -- 
    ack_8903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3290_delayed_13_0_3435_inst_ack_1, ack => sendModule_CP_7983_elements(257)); -- 
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	24 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_Sample/rr
      -- 
    rr_8911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(258), ack => EQ_u3_u1_3447_inst_req_0); -- 
    sendModule_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(24) & sendModule_CP_7983_elements(260);
      gj_sendModule_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: marked-predecessors 
    -- CP-element group 259: 	360 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	261 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_update_start_
      -- CP-element group 259: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_Update/cr
      -- 
    cr_8916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(259), ack => EQ_u3_u1_3447_inst_req_1); -- 
    sendModule_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	22 
    -- CP-element group 260: 	258 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_Sample/ra
      -- 
    ra_8912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3447_inst_ack_0, ack => sendModule_CP_7983_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	259 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	358 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3447_Update/ca
      -- 
    ca_8917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3447_inst_ack_1, ack => sendModule_CP_7983_elements(261)); -- 
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	157 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	264 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_Sample/req
      -- 
    req_8925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(262), ack => W_output_data1_3298_delayed_13_0_3449_inst_req_0); -- 
    sendModule_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(157) & sendModule_CP_7983_elements(264);
      gj_sendModule_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: marked-predecessors 
    -- CP-element group 263: 	360 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	265 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_update_start_
      -- CP-element group 263: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_Update/req
      -- 
    req_8930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(263), ack => W_output_data1_3298_delayed_13_0_3449_inst_req_1); -- 
    sendModule_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: 	155 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_Sample/ack
      -- 
    ack_8926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3298_delayed_13_0_3449_inst_ack_0, ack => sendModule_CP_7983_elements(264)); -- 
    -- CP-element group 265:  transition  input  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	358 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3451_Update/ack
      -- 
    ack_8931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3298_delayed_13_0_3449_inst_ack_1, ack => sendModule_CP_7983_elements(265)); -- 
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	24 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_Sample/rr
      -- 
    rr_8939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(266), ack => EQ_u3_u1_3461_inst_req_0); -- 
    sendModule_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(24) & sendModule_CP_7983_elements(268);
      gj_sendModule_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: marked-predecessors 
    -- CP-element group 267: 	360 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	269 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_update_start_
      -- CP-element group 267: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_Update/cr
      -- 
    cr_8944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(267), ack => EQ_u3_u1_3461_inst_req_1); -- 
    sendModule_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	22 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_Sample/ra
      -- 
    ra_8940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3461_inst_ack_0, ack => sendModule_CP_7983_elements(268)); -- 
    -- CP-element group 269:  transition  input  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	267 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	358 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3461_Update/ca
      -- 
    ca_8945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3461_inst_ack_1, ack => sendModule_CP_7983_elements(269)); -- 
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	157 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	272 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_Sample/req
      -- 
    req_8953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(270), ack => W_output_data1_3306_delayed_13_0_3463_inst_req_0); -- 
    sendModule_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(157) & sendModule_CP_7983_elements(272);
      gj_sendModule_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: marked-predecessors 
    -- CP-element group 271: 	360 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	273 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_update_start_
      -- CP-element group 271: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_Update/req
      -- 
    req_8958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(271), ack => W_output_data1_3306_delayed_13_0_3463_inst_req_1); -- 
    sendModule_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: 	155 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_Sample/ack
      -- 
    ack_8954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3306_delayed_13_0_3463_inst_ack_0, ack => sendModule_CP_7983_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	358 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3465_Update/ack
      -- 
    ack_8959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3306_delayed_13_0_3463_inst_ack_1, ack => sendModule_CP_7983_elements(273)); -- 
    -- CP-element group 274:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	24 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	276 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_Sample/rr
      -- 
    rr_8967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(274), ack => EQ_u3_u1_3475_inst_req_0); -- 
    sendModule_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(24) & sendModule_CP_7983_elements(276);
      gj_sendModule_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: marked-predecessors 
    -- CP-element group 275: 	360 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_update_start_
      -- CP-element group 275: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_Update/cr
      -- 
    cr_8972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(275), ack => EQ_u3_u1_3475_inst_req_1); -- 
    sendModule_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: marked-successors 
    -- CP-element group 276: 	22 
    -- CP-element group 276: 	274 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_sample_completed_
      -- CP-element group 276: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_Sample/ra
      -- 
    ra_8968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3475_inst_ack_0, ack => sendModule_CP_7983_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	358 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_Update/$exit
      -- CP-element group 277: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3475_Update/ca
      -- 
    ca_8973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3475_inst_ack_1, ack => sendModule_CP_7983_elements(277)); -- 
    -- CP-element group 278:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	157 
    -- CP-element group 278: marked-predecessors 
    -- CP-element group 278: 	280 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_Sample/req
      -- 
    req_8981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(278), ack => W_output_data1_3314_delayed_13_0_3477_inst_req_0); -- 
    sendModule_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(157) & sendModule_CP_7983_elements(280);
      gj_sendModule_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: marked-predecessors 
    -- CP-element group 279: 	360 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_update_start_
      -- CP-element group 279: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_Update/req
      -- 
    req_8986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(279), ack => W_output_data1_3314_delayed_13_0_3477_inst_req_1); -- 
    sendModule_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: 	155 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_sample_completed_
      -- CP-element group 280: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_Sample/$exit
      -- CP-element group 280: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_Sample/ack
      -- 
    ack_8982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3314_delayed_13_0_3477_inst_ack_0, ack => sendModule_CP_7983_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	358 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_update_completed_
      -- CP-element group 281: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_Update/$exit
      -- CP-element group 281: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3479_Update/ack
      -- 
    ack_8987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3314_delayed_13_0_3477_inst_ack_1, ack => sendModule_CP_7983_elements(281)); -- 
    -- CP-element group 282:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	24 
    -- CP-element group 282: marked-predecessors 
    -- CP-element group 282: 	284 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_sample_start_
      -- CP-element group 282: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_Sample/rr
      -- 
    rr_8995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(282), ack => EQ_u3_u1_3489_inst_req_0); -- 
    sendModule_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(24) & sendModule_CP_7983_elements(284);
      gj_sendModule_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: marked-predecessors 
    -- CP-element group 283: 	360 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	285 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_update_start_
      -- CP-element group 283: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_Update/cr
      -- 
    cr_9000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(283), ack => EQ_u3_u1_3489_inst_req_1); -- 
    sendModule_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: successors 
    -- CP-element group 284: marked-successors 
    -- CP-element group 284: 	22 
    -- CP-element group 284: 	282 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_Sample/ra
      -- 
    ra_8996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3489_inst_ack_0, ack => sendModule_CP_7983_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	283 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	358 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3489_Update/ca
      -- 
    ca_9001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3489_inst_ack_1, ack => sendModule_CP_7983_elements(285)); -- 
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	157 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	288 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_sample_start_
      -- CP-element group 286: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_Sample/req
      -- 
    req_9009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(286), ack => W_output_data1_3322_delayed_13_0_3491_inst_req_0); -- 
    sendModule_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(157) & sendModule_CP_7983_elements(288);
      gj_sendModule_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: marked-predecessors 
    -- CP-element group 287: 	360 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	289 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_update_start_
      -- CP-element group 287: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_Update/req
      -- 
    req_9014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(287), ack => W_output_data1_3322_delayed_13_0_3491_inst_req_1); -- 
    sendModule_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: 	155 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_Sample/ack
      -- 
    ack_9010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3322_delayed_13_0_3491_inst_ack_0, ack => sendModule_CP_7983_elements(288)); -- 
    -- CP-element group 289:  transition  input  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	287 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	358 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3493_Update/ack
      -- 
    ack_9015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3322_delayed_13_0_3491_inst_ack_1, ack => sendModule_CP_7983_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	43 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_Sample/rr
      -- 
    rr_9023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(290), ack => EQ_u3_u1_3503_inst_req_0); -- 
    sendModule_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(43) & sendModule_CP_7983_elements(292);
      gj_sendModule_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: marked-predecessors 
    -- CP-element group 291: 	372 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_Update/cr
      -- CP-element group 291: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_update_start_
      -- 
    cr_9028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(291), ack => EQ_u3_u1_3503_inst_req_1); -- 
    sendModule_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	39 
    -- CP-element group 292: 	290 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_sample_completed_
      -- CP-element group 292: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_Sample/ra
      -- 
    ra_9024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3503_inst_ack_0, ack => sendModule_CP_7983_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	370 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_Update/ca
      -- CP-element group 293: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3503_update_completed_
      -- 
    ca_9029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3503_inst_ack_1, ack => sendModule_CP_7983_elements(293)); -- 
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	161 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_sample_start_
      -- 
    req_9037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(294), ack => W_output_data2_3330_delayed_13_0_3505_inst_req_0); -- 
    sendModule_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(161) & sendModule_CP_7983_elements(296);
      gj_sendModule_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: marked-predecessors 
    -- CP-element group 295: 	372 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	297 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_Update/req
      -- CP-element group 295: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_update_start_
      -- 
    req_9042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(295), ack => W_output_data2_3330_delayed_13_0_3505_inst_req_1); -- 
    sendModule_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: 	159 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_Sample/ack
      -- CP-element group 296: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_sample_completed_
      -- 
    ack_9038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3330_delayed_13_0_3505_inst_ack_0, ack => sendModule_CP_7983_elements(296)); -- 
    -- CP-element group 297:  transition  input  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	295 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	370 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_Update/ack
      -- CP-element group 297: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3507_update_completed_
      -- 
    ack_9043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3330_delayed_13_0_3505_inst_ack_1, ack => sendModule_CP_7983_elements(297)); -- 
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	43 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_Sample/rr
      -- CP-element group 298: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_Sample/$entry
      -- 
    rr_9051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(298), ack => EQ_u3_u1_3517_inst_req_0); -- 
    sendModule_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(43) & sendModule_CP_7983_elements(300);
      gj_sendModule_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: marked-predecessors 
    -- CP-element group 299: 	372 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	301 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_Update/cr
      -- CP-element group 299: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_update_start_
      -- 
    cr_9056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(299), ack => EQ_u3_u1_3517_inst_req_1); -- 
    sendModule_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	39 
    -- CP-element group 300: 	298 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_Sample/ra
      -- CP-element group 300: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_Sample/$exit
      -- 
    ra_9052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3517_inst_ack_0, ack => sendModule_CP_7983_elements(300)); -- 
    -- CP-element group 301:  transition  input  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	299 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	370 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3517_Update/ca
      -- 
    ca_9057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3517_inst_ack_1, ack => sendModule_CP_7983_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	161 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	304 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_sample_start_
      -- 
    req_9065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(302), ack => W_output_data2_3338_delayed_13_0_3519_inst_req_0); -- 
    sendModule_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(161) & sendModule_CP_7983_elements(304);
      gj_sendModule_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: marked-predecessors 
    -- CP-element group 303: 	372 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	305 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_Update/req
      -- CP-element group 303: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_update_start_
      -- 
    req_9070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(303), ack => W_output_data2_3338_delayed_13_0_3519_inst_req_1); -- 
    sendModule_cp_element_group_303: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_303"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_303 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(303), clk => clk, reset => reset); --
    end block;
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: 	159 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_Sample/$exit
      -- CP-element group 304: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_Sample/ack
      -- CP-element group 304: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_sample_completed_
      -- 
    ack_9066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3338_delayed_13_0_3519_inst_ack_0, ack => sendModule_CP_7983_elements(304)); -- 
    -- CP-element group 305:  transition  input  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	303 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	370 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_update_completed_
      -- CP-element group 305: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_Update/$exit
      -- CP-element group 305: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3521_Update/ack
      -- 
    ack_9071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3338_delayed_13_0_3519_inst_ack_1, ack => sendModule_CP_7983_elements(305)); -- 
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	43 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_Sample/rr
      -- 
    rr_9079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(306), ack => EQ_u3_u1_3531_inst_req_0); -- 
    sendModule_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(43) & sendModule_CP_7983_elements(308);
      gj_sendModule_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: marked-predecessors 
    -- CP-element group 307: 	372 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	309 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_Update/cr
      -- CP-element group 307: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_update_start_
      -- 
    cr_9084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(307), ack => EQ_u3_u1_3531_inst_req_1); -- 
    sendModule_cp_element_group_307: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_307"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_307 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(307), clk => clk, reset => reset); --
    end block;
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	39 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_Sample/ra
      -- CP-element group 308: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_sample_completed_
      -- CP-element group 308: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_Sample/$exit
      -- 
    ra_9080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3531_inst_ack_0, ack => sendModule_CP_7983_elements(308)); -- 
    -- CP-element group 309:  transition  input  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	307 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	370 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_Update/$exit
      -- CP-element group 309: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_Update/ca
      -- CP-element group 309: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3531_update_completed_
      -- 
    ca_9085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3531_inst_ack_1, ack => sendModule_CP_7983_elements(309)); -- 
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	161 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_Sample/$entry
      -- 
    req_9093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(310), ack => W_output_data2_3346_delayed_13_0_3533_inst_req_0); -- 
    sendModule_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(161) & sendModule_CP_7983_elements(312);
      gj_sendModule_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: marked-predecessors 
    -- CP-element group 311: 	372 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	313 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_Update/req
      -- CP-element group 311: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_update_start_
      -- 
    req_9098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(311), ack => W_output_data2_3346_delayed_13_0_3533_inst_req_1); -- 
    sendModule_cp_element_group_311: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_311"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_311 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(311), clk => clk, reset => reset); --
    end block;
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: 	159 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_sample_completed_
      -- CP-element group 312: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_Sample/ack
      -- CP-element group 312: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_Sample/$exit
      -- 
    ack_9094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3346_delayed_13_0_3533_inst_ack_0, ack => sendModule_CP_7983_elements(312)); -- 
    -- CP-element group 313:  transition  input  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	311 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	370 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_Update/ack
      -- CP-element group 313: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3535_update_completed_
      -- 
    ack_9099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3346_delayed_13_0_3533_inst_ack_1, ack => sendModule_CP_7983_elements(313)); -- 
    -- CP-element group 314:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	43 
    -- CP-element group 314: marked-predecessors 
    -- CP-element group 314: 	316 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_Sample/rr
      -- CP-element group 314: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_Sample/$entry
      -- CP-element group 314: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_sample_start_
      -- 
    rr_9107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(314), ack => EQ_u3_u1_3545_inst_req_0); -- 
    sendModule_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(43) & sendModule_CP_7983_elements(316);
      gj_sendModule_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: marked-predecessors 
    -- CP-element group 315: 	372 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_Update/cr
      -- CP-element group 315: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_update_start_
      -- 
    cr_9112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(315), ack => EQ_u3_u1_3545_inst_req_1); -- 
    sendModule_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: successors 
    -- CP-element group 316: marked-successors 
    -- CP-element group 316: 	39 
    -- CP-element group 316: 	314 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_Sample/$exit
      -- CP-element group 316: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_Sample/ra
      -- CP-element group 316: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_sample_completed_
      -- 
    ra_9108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3545_inst_ack_0, ack => sendModule_CP_7983_elements(316)); -- 
    -- CP-element group 317:  transition  input  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	370 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_Update/$exit
      -- CP-element group 317: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_Update/ca
      -- CP-element group 317: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3545_update_completed_
      -- 
    ca_9113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3545_inst_ack_1, ack => sendModule_CP_7983_elements(317)); -- 
    -- CP-element group 318:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	161 
    -- CP-element group 318: marked-predecessors 
    -- CP-element group 318: 	320 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	320 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_sample_start_
      -- CP-element group 318: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_Sample/$entry
      -- CP-element group 318: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_Sample/req
      -- 
    req_9121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(318), ack => W_output_data2_3354_delayed_13_0_3547_inst_req_0); -- 
    sendModule_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(161) & sendModule_CP_7983_elements(320);
      gj_sendModule_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: marked-predecessors 
    -- CP-element group 319: 	372 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_update_start_
      -- CP-element group 319: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_Update/req
      -- 
    req_9126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(319), ack => W_output_data2_3354_delayed_13_0_3547_inst_req_1); -- 
    sendModule_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: successors 
    -- CP-element group 320: marked-successors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: 	159 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_Sample/ack
      -- 
    ack_9122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3354_delayed_13_0_3547_inst_ack_0, ack => sendModule_CP_7983_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	370 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3549_Update/ack
      -- 
    ack_9127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3354_delayed_13_0_3547_inst_ack_1, ack => sendModule_CP_7983_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	43 
    -- CP-element group 322: marked-predecessors 
    -- CP-element group 322: 	324 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_Sample/rr
      -- 
    rr_9135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(322), ack => EQ_u3_u1_3559_inst_req_0); -- 
    sendModule_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(43) & sendModule_CP_7983_elements(324);
      gj_sendModule_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: marked-predecessors 
    -- CP-element group 323: 	372 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_update_start_
      -- CP-element group 323: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_Update/cr
      -- 
    cr_9140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(323), ack => EQ_u3_u1_3559_inst_req_1); -- 
    sendModule_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: successors 
    -- CP-element group 324: marked-successors 
    -- CP-element group 324: 	39 
    -- CP-element group 324: 	322 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_sample_completed_
      -- CP-element group 324: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_Sample/ra
      -- 
    ra_9136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3559_inst_ack_0, ack => sendModule_CP_7983_elements(324)); -- 
    -- CP-element group 325:  transition  input  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	370 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_update_completed_
      -- CP-element group 325: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3559_Update/ca
      -- 
    ca_9141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3559_inst_ack_1, ack => sendModule_CP_7983_elements(325)); -- 
    -- CP-element group 326:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	161 
    -- CP-element group 326: marked-predecessors 
    -- CP-element group 326: 	328 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_Sample/req
      -- 
    req_9149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(326), ack => W_output_data2_3362_delayed_13_0_3561_inst_req_0); -- 
    sendModule_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(161) & sendModule_CP_7983_elements(328);
      gj_sendModule_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: marked-predecessors 
    -- CP-element group 327: 	372 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	329 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_update_start_
      -- CP-element group 327: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_Update/req
      -- 
    req_9154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(327), ack => W_output_data2_3362_delayed_13_0_3561_inst_req_1); -- 
    sendModule_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: successors 
    -- CP-element group 328: marked-successors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: 	159 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_sample_completed_
      -- CP-element group 328: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_Sample/$exit
      -- CP-element group 328: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_Sample/ack
      -- 
    ack_9150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3362_delayed_13_0_3561_inst_ack_0, ack => sendModule_CP_7983_elements(328)); -- 
    -- CP-element group 329:  transition  input  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	327 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	370 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_update_completed_
      -- CP-element group 329: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_Update/$exit
      -- CP-element group 329: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3563_Update/ack
      -- 
    ack_9155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3362_delayed_13_0_3561_inst_ack_1, ack => sendModule_CP_7983_elements(329)); -- 
    -- CP-element group 330:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	43 
    -- CP-element group 330: marked-predecessors 
    -- CP-element group 330: 	332 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	332 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_sample_start_
      -- CP-element group 330: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_Sample/rr
      -- CP-element group 330: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_Sample/$entry
      -- 
    rr_9163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(330), ack => EQ_u3_u1_3573_inst_req_0); -- 
    sendModule_cp_element_group_330: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_330"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(43) & sendModule_CP_7983_elements(332);
      gj_sendModule_cp_element_group_330 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(330), clk => clk, reset => reset); --
    end block;
    -- CP-element group 331:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: marked-predecessors 
    -- CP-element group 331: 	372 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	333 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_Update/cr
      -- CP-element group 331: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_update_start_
      -- 
    cr_9168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(331), ack => EQ_u3_u1_3573_inst_req_1); -- 
    sendModule_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: successors 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	39 
    -- CP-element group 332: 	330 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_sample_completed_
      -- CP-element group 332: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_Sample/ra
      -- CP-element group 332: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_Sample/$exit
      -- 
    ra_9164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3573_inst_ack_0, ack => sendModule_CP_7983_elements(332)); -- 
    -- CP-element group 333:  transition  input  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	331 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	370 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_Update/$exit
      -- CP-element group 333: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_Update/ca
      -- CP-element group 333: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3573_update_completed_
      -- 
    ca_9169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3573_inst_ack_1, ack => sendModule_CP_7983_elements(333)); -- 
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	161 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_Sample/req
      -- CP-element group 334: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_Sample/$entry
      -- 
    req_9177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(334), ack => W_output_data2_3370_delayed_13_0_3575_inst_req_0); -- 
    sendModule_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(161) & sendModule_CP_7983_elements(336);
      gj_sendModule_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: marked-predecessors 
    -- CP-element group 335: 	372 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_Update/req
      -- CP-element group 335: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_update_start_
      -- 
    req_9182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(335), ack => W_output_data2_3370_delayed_13_0_3575_inst_req_1); -- 
    sendModule_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: 	159 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_sample_completed_
      -- CP-element group 336: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_Sample/ack
      -- CP-element group 336: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_Sample/$exit
      -- 
    ack_9178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3370_delayed_13_0_3575_inst_ack_0, ack => sendModule_CP_7983_elements(336)); -- 
    -- CP-element group 337:  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	370 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_Update/ack
      -- CP-element group 337: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_Update/$exit
      -- CP-element group 337: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3577_update_completed_
      -- 
    ack_9183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3370_delayed_13_0_3575_inst_ack_1, ack => sendModule_CP_7983_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	43 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_Sample/rr
      -- CP-element group 338: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_sample_start_
      -- 
    rr_9191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(338), ack => EQ_u3_u1_3587_inst_req_0); -- 
    sendModule_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(43) & sendModule_CP_7983_elements(340);
      gj_sendModule_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	372 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_Update/cr
      -- CP-element group 339: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_update_start_
      -- 
    cr_9196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(339), ack => EQ_u3_u1_3587_inst_req_1); -- 
    sendModule_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	39 
    -- CP-element group 340: 	338 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_Sample/ra
      -- CP-element group 340: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_sample_completed_
      -- 
    ra_9192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3587_inst_ack_0, ack => sendModule_CP_7983_elements(340)); -- 
    -- CP-element group 341:  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	370 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_Update/ca
      -- CP-element group 341: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3587_update_completed_
      -- 
    ca_9197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3587_inst_ack_1, ack => sendModule_CP_7983_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	161 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_Sample/req
      -- CP-element group 342: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_sample_start_
      -- 
    req_9205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(342), ack => W_output_data2_3378_delayed_13_0_3589_inst_req_0); -- 
    sendModule_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(161) & sendModule_CP_7983_elements(344);
      gj_sendModule_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	372 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_Update/req
      -- CP-element group 343: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_update_start_
      -- 
    req_9210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(343), ack => W_output_data2_3378_delayed_13_0_3589_inst_req_1); -- 
    sendModule_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: 	159 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_Sample/ack
      -- CP-element group 344: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_Sample/$exit
      -- CP-element group 344: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_sample_completed_
      -- 
    ack_9206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3378_delayed_13_0_3589_inst_ack_0, ack => sendModule_CP_7983_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	370 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_Update/$exit
      -- CP-element group 345: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_Update/ack
      -- CP-element group 345: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3591_update_completed_
      -- 
    ack_9211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3378_delayed_13_0_3589_inst_ack_1, ack => sendModule_CP_7983_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	43 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	348 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_Sample/rr
      -- 
    rr_9219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(346), ack => EQ_u3_u1_3601_inst_req_0); -- 
    sendModule_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(43) & sendModule_CP_7983_elements(348);
      gj_sendModule_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: marked-predecessors 
    -- CP-element group 347: 	372 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	349 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_update_start_
      -- CP-element group 347: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_Update/cr
      -- CP-element group 347: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_Update/$entry
      -- 
    cr_9224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(347), ack => EQ_u3_u1_3601_inst_req_1); -- 
    sendModule_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: successors 
    -- CP-element group 348: marked-successors 
    -- CP-element group 348: 	39 
    -- CP-element group 348: 	346 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_sample_completed_
      -- CP-element group 348: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_Sample/$exit
      -- CP-element group 348: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_Sample/ra
      -- 
    ra_9220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3601_inst_ack_0, ack => sendModule_CP_7983_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	347 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	370 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_update_completed_
      -- CP-element group 349: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_Update/ca
      -- CP-element group 349: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/EQ_u3_u1_3601_Update/$exit
      -- 
    ca_9225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3601_inst_ack_1, ack => sendModule_CP_7983_elements(349)); -- 
    -- CP-element group 350:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	161 
    -- CP-element group 350: marked-predecessors 
    -- CP-element group 350: 	352 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_Sample/req
      -- CP-element group 350: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_Sample/$entry
      -- CP-element group 350: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_sample_start_
      -- 
    req_9233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(350), ack => W_output_data2_3386_delayed_13_0_3603_inst_req_0); -- 
    sendModule_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(161) & sendModule_CP_7983_elements(352);
      gj_sendModule_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: marked-predecessors 
    -- CP-element group 351: 	372 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_Update/req
      -- CP-element group 351: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_Update/$entry
      -- CP-element group 351: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_update_start_
      -- 
    req_9238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(351), ack => W_output_data2_3386_delayed_13_0_3603_inst_req_1); -- 
    sendModule_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: successors 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: 	159 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_sample_completed_
      -- 
    ack_9234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3386_delayed_13_0_3603_inst_ack_0, ack => sendModule_CP_7983_elements(352)); -- 
    -- CP-element group 353:  transition  input  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	370 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_Update/ack
      -- CP-element group 353: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3605_update_completed_
      -- 
    ack_9239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3386_delayed_13_0_3603_inst_ack_1, ack => sendModule_CP_7983_elements(353)); -- 
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	134 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_Sample/$entry
      -- CP-element group 354: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_Sample/req
      -- CP-element group 354: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_sample_start_
      -- 
    req_9247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(354), ack => W_fetch_addr1_3390_delayed_8_0_3612_inst_req_0); -- 
    sendModule_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(134) & sendModule_CP_7983_elements(356);
      gj_sendModule_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: marked-predecessors 
    -- CP-element group 355: 	364 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	357 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_Update/req
      -- CP-element group 355: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_update_start_
      -- 
    req_9252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(355), ack => W_fetch_addr1_3390_delayed_8_0_3612_inst_req_1); -- 
    sendModule_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(364);
      gj_sendModule_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: 	129 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_Sample/ack
      -- CP-element group 356: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_sample_completed_
      -- 
    ack_9248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr1_3390_delayed_8_0_3612_inst_ack_0, ack => sendModule_CP_7983_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	355 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	362 
    -- CP-element group 357:  members (19) 
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_base_addr_resize/base_resize_ack
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_base_plus_offset/$entry
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_base_plus_offset/$exit
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_base_plus_offset/sum_rename_req
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_base_plus_offset/sum_rename_ack
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3614_Update/ack
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_word_addrgen/$entry
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_word_addrgen/$exit
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_word_addrgen/root_register_req
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_base_addr_resize/base_resize_req
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_base_addr_resize/$exit
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_base_addr_resize/$entry
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_base_address_resized
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_root_address_calculated
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_word_address_calculated
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_base_address_calculated
      -- CP-element group 357: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_word_addrgen/root_register_ack
      -- 
    ack_9253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr1_3390_delayed_8_0_3612_inst_ack_1, ack => sendModule_CP_7983_elements(357)); -- 
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	165 
    -- CP-element group 358: 	169 
    -- CP-element group 358: 	173 
    -- CP-element group 358: 	177 
    -- CP-element group 358: 	269 
    -- CP-element group 358: 	273 
    -- CP-element group 358: 	277 
    -- CP-element group 358: 	281 
    -- CP-element group 358: 	285 
    -- CP-element group 358: 	289 
    -- CP-element group 358: 	253 
    -- CP-element group 358: 	257 
    -- CP-element group 358: 	261 
    -- CP-element group 358: 	265 
    -- CP-element group 358: 	233 
    -- CP-element group 358: 	237 
    -- CP-element group 358: 	241 
    -- CP-element group 358: 	245 
    -- CP-element group 358: 	249 
    -- CP-element group 358: 	181 
    -- CP-element group 358: 	185 
    -- CP-element group 358: 	189 
    -- CP-element group 358: 	193 
    -- CP-element group 358: 	229 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_Sample/rr
      -- 
    rr_9261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(358), ack => CONCAT_u32_u64_3631_inst_req_0); -- 
    sendModule_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 24) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1);
      constant place_markings: IntegerArray(0 to 24)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 1);
      constant place_delays: IntegerArray(0 to 24) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 25); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(165) & sendModule_CP_7983_elements(169) & sendModule_CP_7983_elements(173) & sendModule_CP_7983_elements(177) & sendModule_CP_7983_elements(269) & sendModule_CP_7983_elements(273) & sendModule_CP_7983_elements(277) & sendModule_CP_7983_elements(281) & sendModule_CP_7983_elements(285) & sendModule_CP_7983_elements(289) & sendModule_CP_7983_elements(253) & sendModule_CP_7983_elements(257) & sendModule_CP_7983_elements(261) & sendModule_CP_7983_elements(265) & sendModule_CP_7983_elements(233) & sendModule_CP_7983_elements(237) & sendModule_CP_7983_elements(241) & sendModule_CP_7983_elements(245) & sendModule_CP_7983_elements(249) & sendModule_CP_7983_elements(181) & sendModule_CP_7983_elements(185) & sendModule_CP_7983_elements(189) & sendModule_CP_7983_elements(193) & sendModule_CP_7983_elements(229) & sendModule_CP_7983_elements(360);
      gj_sendModule_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 25, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: marked-predecessors 
    -- CP-element group 359: 	364 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_update_start_
      -- CP-element group 359: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_Update/cr
      -- 
    cr_9266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(359), ack => CONCAT_u32_u64_3631_inst_req_1); -- 
    sendModule_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(364);
      gj_sendModule_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	167 
    -- CP-element group 360: 	171 
    -- CP-element group 360: 	175 
    -- CP-element group 360: 	271 
    -- CP-element group 360: 	275 
    -- CP-element group 360: 	279 
    -- CP-element group 360: 	283 
    -- CP-element group 360: 	287 
    -- CP-element group 360: 	251 
    -- CP-element group 360: 	255 
    -- CP-element group 360: 	259 
    -- CP-element group 360: 	263 
    -- CP-element group 360: 	267 
    -- CP-element group 360: 	358 
    -- CP-element group 360: 	235 
    -- CP-element group 360: 	239 
    -- CP-element group 360: 	243 
    -- CP-element group 360: 	247 
    -- CP-element group 360: 	179 
    -- CP-element group 360: 	183 
    -- CP-element group 360: 	187 
    -- CP-element group 360: 	191 
    -- CP-element group 360: 	227 
    -- CP-element group 360: 	231 
    -- CP-element group 360: 	163 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_Sample/ra
      -- CP-element group 360: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_sample_completed_
      -- CP-element group 360: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_Sample/$exit
      -- 
    ra_9262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3631_inst_ack_0, ack => sendModule_CP_7983_elements(360)); -- 
    -- CP-element group 361:  transition  input  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_update_completed_
      -- CP-element group 361: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3631_Update/ca
      -- 
    ca_9267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3631_inst_ack_1, ack => sendModule_CP_7983_elements(361)); -- 
    -- CP-element group 362:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	383 
    -- CP-element group 362: 	384 
    -- CP-element group 362: 	357 
    -- CP-element group 362: 	361 
    -- CP-element group 362: marked-predecessors 
    -- CP-element group 362: 	364 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (9) 
      -- CP-element group 362: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/word_access_start/word_0/rr
      -- CP-element group 362: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/word_access_start/word_0/$entry
      -- CP-element group 362: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/word_access_start/$entry
      -- CP-element group 362: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/ptr_deref_3616_Split/split_ack
      -- CP-element group 362: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/ptr_deref_3616_Split/split_req
      -- CP-element group 362: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/ptr_deref_3616_Split/$exit
      -- CP-element group 362: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/ptr_deref_3616_Split/$entry
      -- CP-element group 362: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/$entry
      -- 
    rr_9305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(362), ack => ptr_deref_3616_store_0_req_0); -- 
    sendModule_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(383) & sendModule_CP_7983_elements(384) & sendModule_CP_7983_elements(357) & sendModule_CP_7983_elements(361) & sendModule_CP_7983_elements(364);
      gj_sendModule_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: marked-predecessors 
    -- CP-element group 363: 	365 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	365 
    -- CP-element group 363:  members (5) 
      -- CP-element group 363: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Update/word_access_complete/word_0/cr
      -- CP-element group 363: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Update/word_access_complete/word_0/$entry
      -- CP-element group 363: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Update/word_access_complete/$entry
      -- CP-element group 363: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_update_start_
      -- 
    cr_9316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(363), ack => ptr_deref_3616_store_0_req_1); -- 
    sendModule_cp_element_group_363: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_363"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(365);
      gj_sendModule_cp_element_group_363 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 364:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	385 
    -- CP-element group 364: marked-successors 
    -- CP-element group 364: 	355 
    -- CP-element group 364: 	359 
    -- CP-element group 364: 	362 
    -- CP-element group 364:  members (5) 
      -- CP-element group 364: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/word_access_start/word_0/ra
      -- CP-element group 364: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/word_access_start/word_0/$exit
      -- CP-element group 364: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/word_access_start/$exit
      -- CP-element group 364: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_sample_completed_
      -- CP-element group 364: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Sample/$exit
      -- 
    ra_9306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3616_store_0_ack_0, ack => sendModule_CP_7983_elements(364)); -- 
    -- CP-element group 365:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	363 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	386 
    -- CP-element group 365: marked-successors 
    -- CP-element group 365: 	363 
    -- CP-element group 365:  members (5) 
      -- CP-element group 365: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Update/word_access_complete/word_0/ca
      -- CP-element group 365: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Update/word_access_complete/word_0/$exit
      -- CP-element group 365: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Update/word_access_complete/$exit
      -- CP-element group 365: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_update_completed_
      -- 
    ca_9317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3616_store_0_ack_1, ack => sendModule_CP_7983_elements(365)); -- 
    -- CP-element group 366:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	141 
    -- CP-element group 366: marked-predecessors 
    -- CP-element group 366: 	368 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	368 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_Sample/req
      -- CP-element group 366: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_sample_start_
      -- 
    req_9325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(366), ack => W_fetch_addr2_3408_delayed_8_0_3633_inst_req_0); -- 
    sendModule_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(141) & sendModule_CP_7983_elements(368);
      gj_sendModule_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	376 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_Update/req
      -- CP-element group 367: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_update_start_
      -- 
    req_9330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(367), ack => W_fetch_addr2_3408_delayed_8_0_3633_inst_req_1); -- 
    sendModule_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(376);
      gj_sendModule_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: successors 
    -- CP-element group 368: marked-successors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: 	136 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_Sample/ack
      -- CP-element group 368: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_sample_completed_
      -- 
    ack_9326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr2_3408_delayed_8_0_3633_inst_ack_0, ack => sendModule_CP_7983_elements(368)); -- 
    -- CP-element group 369:  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	374 
    -- CP-element group 369:  members (19) 
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_Update/ack
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_base_address_resized
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_word_addrgen/root_register_req
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_word_addrgen/root_register_ack
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_word_address_calculated
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_word_addrgen/$entry
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_base_address_calculated
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/assign_stmt_3635_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_base_plus_offset/sum_rename_ack
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_base_plus_offset/sum_rename_req
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_base_plus_offset/$exit
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_base_plus_offset/$entry
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_base_addr_resize/base_resize_ack
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_base_addr_resize/base_resize_req
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_base_addr_resize/$exit
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_base_addr_resize/$entry
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_root_address_calculated
      -- CP-element group 369: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_word_addrgen/$exit
      -- 
    ack_9331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr2_3408_delayed_8_0_3633_inst_ack_1, ack => sendModule_CP_7983_elements(369)); -- 
    -- CP-element group 370:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	293 
    -- CP-element group 370: 	297 
    -- CP-element group 370: 	301 
    -- CP-element group 370: 	305 
    -- CP-element group 370: 	309 
    -- CP-element group 370: 	313 
    -- CP-element group 370: 	317 
    -- CP-element group 370: 	321 
    -- CP-element group 370: 	341 
    -- CP-element group 370: 	345 
    -- CP-element group 370: 	349 
    -- CP-element group 370: 	353 
    -- CP-element group 370: 	325 
    -- CP-element group 370: 	329 
    -- CP-element group 370: 	333 
    -- CP-element group 370: 	337 
    -- CP-element group 370: 	197 
    -- CP-element group 370: 	201 
    -- CP-element group 370: 	205 
    -- CP-element group 370: 	209 
    -- CP-element group 370: 	213 
    -- CP-element group 370: 	217 
    -- CP-element group 370: 	221 
    -- CP-element group 370: 	225 
    -- CP-element group 370: marked-predecessors 
    -- CP-element group 370: 	372 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	372 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_sample_start_
      -- CP-element group 370: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_Sample/$entry
      -- CP-element group 370: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_Sample/rr
      -- 
    rr_9339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(370), ack => CONCAT_u32_u64_3652_inst_req_0); -- 
    sendModule_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 24) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1);
      constant place_markings: IntegerArray(0 to 24)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 1);
      constant place_delays: IntegerArray(0 to 24) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 25); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(293) & sendModule_CP_7983_elements(297) & sendModule_CP_7983_elements(301) & sendModule_CP_7983_elements(305) & sendModule_CP_7983_elements(309) & sendModule_CP_7983_elements(313) & sendModule_CP_7983_elements(317) & sendModule_CP_7983_elements(321) & sendModule_CP_7983_elements(341) & sendModule_CP_7983_elements(345) & sendModule_CP_7983_elements(349) & sendModule_CP_7983_elements(353) & sendModule_CP_7983_elements(325) & sendModule_CP_7983_elements(329) & sendModule_CP_7983_elements(333) & sendModule_CP_7983_elements(337) & sendModule_CP_7983_elements(197) & sendModule_CP_7983_elements(201) & sendModule_CP_7983_elements(205) & sendModule_CP_7983_elements(209) & sendModule_CP_7983_elements(213) & sendModule_CP_7983_elements(217) & sendModule_CP_7983_elements(221) & sendModule_CP_7983_elements(225) & sendModule_CP_7983_elements(372);
      gj_sendModule_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 25, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: marked-predecessors 
    -- CP-element group 371: 	376 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	373 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_update_start_
      -- CP-element group 371: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_Update/cr
      -- CP-element group 371: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_Update/$entry
      -- 
    cr_9344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(371), ack => CONCAT_u32_u64_3652_inst_req_1); -- 
    sendModule_cp_element_group_371: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_371"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(376);
      gj_sendModule_cp_element_group_371 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(371), clk => clk, reset => reset); --
    end block;
    -- CP-element group 372:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	370 
    -- CP-element group 372: successors 
    -- CP-element group 372: marked-successors 
    -- CP-element group 372: 	370 
    -- CP-element group 372: 	291 
    -- CP-element group 372: 	295 
    -- CP-element group 372: 	299 
    -- CP-element group 372: 	303 
    -- CP-element group 372: 	307 
    -- CP-element group 372: 	311 
    -- CP-element group 372: 	315 
    -- CP-element group 372: 	319 
    -- CP-element group 372: 	343 
    -- CP-element group 372: 	347 
    -- CP-element group 372: 	351 
    -- CP-element group 372: 	323 
    -- CP-element group 372: 	327 
    -- CP-element group 372: 	331 
    -- CP-element group 372: 	335 
    -- CP-element group 372: 	339 
    -- CP-element group 372: 	195 
    -- CP-element group 372: 	199 
    -- CP-element group 372: 	203 
    -- CP-element group 372: 	207 
    -- CP-element group 372: 	211 
    -- CP-element group 372: 	215 
    -- CP-element group 372: 	219 
    -- CP-element group 372: 	223 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_Sample/ra
      -- 
    ra_9340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3652_inst_ack_0, ack => sendModule_CP_7983_elements(372)); -- 
    -- CP-element group 373:  transition  input  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	371 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_Update/ca
      -- CP-element group 373: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/CONCAT_u32_u64_3652_Update/$exit
      -- 
    ca_9345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3652_inst_ack_1, ack => sendModule_CP_7983_elements(373)); -- 
    -- CP-element group 374:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	369 
    -- CP-element group 374: 	373 
    -- CP-element group 374: 	385 
    -- CP-element group 374: marked-predecessors 
    -- CP-element group 374: 	376 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	376 
    -- CP-element group 374:  members (9) 
      -- CP-element group 374: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/ptr_deref_3637_Split/$entry
      -- CP-element group 374: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/ptr_deref_3637_Split/$exit
      -- CP-element group 374: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/ptr_deref_3637_Split/split_req
      -- CP-element group 374: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/ptr_deref_3637_Split/split_ack
      -- CP-element group 374: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/word_access_start/$entry
      -- CP-element group 374: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/word_access_start/word_0/$entry
      -- CP-element group 374: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/word_access_start/word_0/rr
      -- 
    rr_9383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(374), ack => ptr_deref_3637_store_0_req_0); -- 
    sendModule_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(369) & sendModule_CP_7983_elements(373) & sendModule_CP_7983_elements(385) & sendModule_CP_7983_elements(376);
      gj_sendModule_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: marked-predecessors 
    -- CP-element group 375: 	377 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (5) 
      -- CP-element group 375: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_update_start_
      -- CP-element group 375: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Update/word_access_complete/$entry
      -- CP-element group 375: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Update/word_access_complete/word_0/$entry
      -- CP-element group 375: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Update/word_access_complete/word_0/cr
      -- 
    cr_9394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(375), ack => ptr_deref_3637_store_0_req_1); -- 
    sendModule_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(377);
      gj_sendModule_cp_element_group_375 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	374 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	386 
    -- CP-element group 376: marked-successors 
    -- CP-element group 376: 	142 
    -- CP-element group 376: 	367 
    -- CP-element group 376: 	371 
    -- CP-element group 376: 	374 
    -- CP-element group 376: 	146 
    -- CP-element group 376:  members (6) 
      -- CP-element group 376: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/word_access_start/$exit
      -- CP-element group 376: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/word_access_start/word_0/$exit
      -- CP-element group 376: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Sample/word_access_start/word_0/ra
      -- CP-element group 376: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ring_reenable_memory_space_0
      -- 
    ra_9384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3637_store_0_ack_0, ack => sendModule_CP_7983_elements(376)); -- 
    -- CP-element group 377:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	386 
    -- CP-element group 377: marked-successors 
    -- CP-element group 377: 	375 
    -- CP-element group 377:  members (5) 
      -- CP-element group 377: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Update/word_access_complete/$exit
      -- CP-element group 377: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Update/word_access_complete/word_0/$exit
      -- CP-element group 377: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3637_Update/word_access_complete/word_0/ca
      -- 
    ca_9395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3637_store_0_ack_1, ack => sendModule_CP_7983_elements(377)); -- 
    -- CP-element group 378:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	15 
    -- CP-element group 378: marked-predecessors 
    -- CP-element group 378: 	380 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	380 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_Sample/rr
      -- 
    rr_9403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(378), ack => SUB_u16_u16_3657_inst_req_0); -- 
    sendModule_cp_element_group_378: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_378"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(15) & sendModule_CP_7983_elements(380);
      gj_sendModule_cp_element_group_378 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(378), clk => clk, reset => reset); --
    end block;
    -- CP-element group 379:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: marked-predecessors 
    -- CP-element group 379: 	381 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	381 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_update_start_
      -- CP-element group 379: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_Update/cr
      -- 
    cr_9408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(379), ack => SUB_u16_u16_3657_inst_req_1); -- 
    sendModule_cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_379"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7983_elements(381);
      gj_sendModule_cp_element_group_379 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(379), clk => clk, reset => reset); --
    end block;
    -- CP-element group 380:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	378 
    -- CP-element group 380: successors 
    -- CP-element group 380: marked-successors 
    -- CP-element group 380: 	378 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_Sample/ra
      -- 
    ra_9404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3657_inst_ack_0, ack => sendModule_CP_7983_elements(380)); -- 
    -- CP-element group 381:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	379 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	16 
    -- CP-element group 381: marked-successors 
    -- CP-element group 381: 	379 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/SUB_u16_u16_3657_Update/ca
      -- 
    ca_9409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3657_inst_ack_1, ack => sendModule_CP_7983_elements(381)); -- 
    -- CP-element group 382:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	15 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	16 
    -- CP-element group 382:  members (1) 
      -- CP-element group 382: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group sendModule_CP_7983_elements(382) is a control-delay.
    cp_element_382_delay: control_delay_element  generic map(name => " 382_delay", delay_value => 1)  port map(req => sendModule_CP_7983_elements(15), ack => sendModule_CP_7983_elements(382), clk => clk, reset =>reset);
    -- CP-element group 383:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	144 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	362 
    -- CP-element group 383:  members (1) 
      -- CP-element group 383: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3299_ptr_deref_3616_delay
      -- 
    -- Element group sendModule_CP_7983_elements(383) is a control-delay.
    cp_element_383_delay: control_delay_element  generic map(name => " 383_delay", delay_value => 1)  port map(req => sendModule_CP_7983_elements(144), ack => sendModule_CP_7983_elements(383), clk => clk, reset =>reset);
    -- CP-element group 384:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	148 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	362 
    -- CP-element group 384:  members (1) 
      -- CP-element group 384: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3303_ptr_deref_3616_delay
      -- 
    -- Element group sendModule_CP_7983_elements(384) is a control-delay.
    cp_element_384_delay: control_delay_element  generic map(name => " 384_delay", delay_value => 1)  port map(req => sendModule_CP_7983_elements(148), ack => sendModule_CP_7983_elements(384), clk => clk, reset =>reset);
    -- CP-element group 385:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	364 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	374 
    -- CP-element group 385:  members (1) 
      -- CP-element group 385: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/ptr_deref_3616_ptr_deref_3637_delay
      -- 
    -- Element group sendModule_CP_7983_elements(385) is a control-delay.
    cp_element_385_delay: control_delay_element  generic map(name => " 385_delay", delay_value => 1)  port map(req => sendModule_CP_7983_elements(364), ack => sendModule_CP_7983_elements(385), clk => clk, reset =>reset);
    -- CP-element group 386:  join  transition  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	18 
    -- CP-element group 386: 	138 
    -- CP-element group 386: 	376 
    -- CP-element group 386: 	377 
    -- CP-element group 386: 	365 
    -- CP-element group 386: 	123 
    -- CP-element group 386: 	127 
    -- CP-element group 386: 	131 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	12 
    -- CP-element group 386:  members (1) 
      -- CP-element group 386: 	 branch_block_stmt_3145/do_while_stmt_3161/do_while_stmt_3161_loop_body/$exit
      -- 
    sendModule_cp_element_group_386: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_386"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_7983_elements(18) & sendModule_CP_7983_elements(138) & sendModule_CP_7983_elements(376) & sendModule_CP_7983_elements(377) & sendModule_CP_7983_elements(365) & sendModule_CP_7983_elements(123) & sendModule_CP_7983_elements(127) & sendModule_CP_7983_elements(131);
      gj_sendModule_cp_element_group_386 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7983_elements(386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 387:  transition  input  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	11 
    -- CP-element group 387: successors 
    -- CP-element group 387:  members (2) 
      -- CP-element group 387: 	 branch_block_stmt_3145/do_while_stmt_3161/loop_exit/$exit
      -- CP-element group 387: 	 branch_block_stmt_3145/do_while_stmt_3161/loop_exit/ack
      -- 
    ack_9418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3161_branch_ack_0, ack => sendModule_CP_7983_elements(387)); -- 
    -- CP-element group 388:  transition  input  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	11 
    -- CP-element group 388: successors 
    -- CP-element group 388:  members (2) 
      -- CP-element group 388: 	 branch_block_stmt_3145/do_while_stmt_3161/loop_taken/$exit
      -- CP-element group 388: 	 branch_block_stmt_3145/do_while_stmt_3161/loop_taken/ack
      -- 
    ack_9422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3161_branch_ack_1, ack => sendModule_CP_7983_elements(388)); -- 
    -- CP-element group 389:  transition  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	9 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	1 
    -- CP-element group 389:  members (1) 
      -- CP-element group 389: 	 branch_block_stmt_3145/do_while_stmt_3161/$exit
      -- 
    sendModule_CP_7983_elements(389) <= sendModule_CP_7983_elements(9);
    -- CP-element group 390:  transition  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	1 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (6) 
      -- CP-element group 390: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_update_start_
      -- CP-element group 390: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_Sample/ack
      -- CP-element group 390: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_Update/req
      -- 
    ack_9435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3669_inst_ack_0, ack => sendModule_CP_7983_elements(390)); -- 
    req_9439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7983_elements(390), ack => WPIPE_input_done_pipe_3669_inst_req_1); -- 
    -- CP-element group 391:  transition  place  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391:  members (8) 
      -- CP-element group 391: 	 $exit
      -- CP-element group 391: 	 branch_block_stmt_3145/$exit
      -- CP-element group 391: 	 branch_block_stmt_3145/branch_block_stmt_3145__exit__
      -- CP-element group 391: 	 branch_block_stmt_3145/assign_stmt_3671__exit__
      -- CP-element group 391: 	 branch_block_stmt_3145/assign_stmt_3671/$exit
      -- CP-element group 391: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_3145/assign_stmt_3671/WPIPE_input_done_pipe_3669_Update/ack
      -- 
    ack_9440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3669_inst_ack_1, ack => sendModule_CP_7983_elements(391)); -- 
    sendModule_do_while_stmt_3161_terminator_9423: loop_terminator -- 
      generic map (name => " sendModule_do_while_stmt_3161_terminator_9423", max_iterations_in_flight =>15) 
      port map(loop_body_exit => sendModule_CP_7983_elements(12),loop_continue => sendModule_CP_7983_elements(388),loop_terminate => sendModule_CP_7983_elements(387),loop_back => sendModule_CP_7983_elements(10),loop_exit => sendModule_CP_7983_elements(9),clk => clk, reset => reset); -- 
    phi_stmt_3163_phi_seq_8105_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7983_elements(27);
      sendModule_CP_7983_elements(30)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7983_elements(30);
      sendModule_CP_7983_elements(31)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7983_elements(32);
      sendModule_CP_7983_elements(28) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7983_elements(25);
      sendModule_CP_7983_elements(34)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7983_elements(36);
      sendModule_CP_7983_elements(35)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7983_elements(37);
      sendModule_CP_7983_elements(26) <= phi_mux_reqs(1);
      phi_stmt_3163_phi_seq_8105 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3163_phi_seq_8105") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7983_elements(17), 
          phi_sample_ack => sendModule_CP_7983_elements(23), 
          phi_update_req => sendModule_CP_7983_elements(19), 
          phi_update_ack => sendModule_CP_7983_elements(24), 
          phi_mux_ack => sendModule_CP_7983_elements(29), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3168_phi_seq_8159_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7983_elements(46);
      sendModule_CP_7983_elements(49)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7983_elements(53);
      sendModule_CP_7983_elements(50)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7983_elements(54);
      sendModule_CP_7983_elements(47) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7983_elements(44);
      sendModule_CP_7983_elements(55)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7983_elements(57);
      sendModule_CP_7983_elements(56)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7983_elements(58);
      sendModule_CP_7983_elements(45) <= phi_mux_reqs(1);
      phi_stmt_3168_phi_seq_8159 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3168_phi_seq_8159") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7983_elements(40), 
          phi_sample_ack => sendModule_CP_7983_elements(41), 
          phi_update_req => sendModule_CP_7983_elements(42), 
          phi_update_ack => sendModule_CP_7983_elements(43), 
          phi_mux_ack => sendModule_CP_7983_elements(48), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3173_phi_seq_8203_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7983_elements(67);
      sendModule_CP_7983_elements(70)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7983_elements(70);
      sendModule_CP_7983_elements(71)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7983_elements(72);
      sendModule_CP_7983_elements(68) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7983_elements(65);
      sendModule_CP_7983_elements(74)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7983_elements(76);
      sendModule_CP_7983_elements(75)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7983_elements(77);
      sendModule_CP_7983_elements(66) <= phi_mux_reqs(1);
      phi_stmt_3173_phi_seq_8203 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3173_phi_seq_8203") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7983_elements(61), 
          phi_sample_ack => sendModule_CP_7983_elements(62), 
          phi_update_req => sendModule_CP_7983_elements(63), 
          phi_update_ack => sendModule_CP_7983_elements(64), 
          phi_mux_ack => sendModule_CP_7983_elements(69), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3178_phi_seq_8247_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7983_elements(86);
      sendModule_CP_7983_elements(89)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7983_elements(89);
      sendModule_CP_7983_elements(90)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7983_elements(91);
      sendModule_CP_7983_elements(87) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7983_elements(84);
      sendModule_CP_7983_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7983_elements(95);
      sendModule_CP_7983_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7983_elements(96);
      sendModule_CP_7983_elements(85) <= phi_mux_reqs(1);
      phi_stmt_3178_phi_seq_8247 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3178_phi_seq_8247") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7983_elements(80), 
          phi_sample_ack => sendModule_CP_7983_elements(81), 
          phi_update_req => sendModule_CP_7983_elements(82), 
          phi_update_ack => sendModule_CP_7983_elements(83), 
          phi_mux_ack => sendModule_CP_7983_elements(88), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3183_phi_seq_8291_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7983_elements(105);
      sendModule_CP_7983_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7983_elements(108);
      sendModule_CP_7983_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7983_elements(110);
      sendModule_CP_7983_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7983_elements(103);
      sendModule_CP_7983_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7983_elements(114);
      sendModule_CP_7983_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7983_elements(115);
      sendModule_CP_7983_elements(104) <= phi_mux_reqs(1);
      phi_stmt_3183_phi_seq_8291 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3183_phi_seq_8291") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7983_elements(99), 
          phi_sample_ack => sendModule_CP_7983_elements(100), 
          phi_update_req => sendModule_CP_7983_elements(101), 
          phi_update_ack => sendModule_CP_7983_elements(102), 
          phi_mux_ack => sendModule_CP_7983_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_8057_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= sendModule_CP_7983_elements(13);
        preds(1)  <= sendModule_CP_7983_elements(14);
        entry_tmerge_8057 : transition_merge -- 
          generic map(name => " entry_tmerge_8057")
          port map (preds => preds, symbol_out => sendModule_CP_7983_elements(15));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_3211_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3220_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3229_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_3258_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_3268_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_3272_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3623_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3630_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3644_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3651_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_3631_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_3652_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u8_u16_3619_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3622_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3626_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3629_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3640_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3643_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3647_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3650_wire : std_logic_vector(15 downto 0);
    signal EQ_u3_u1_3265_3265_delayed_14_0_3392 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3273_3273_delayed_14_0_3406 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3281_3281_delayed_14_0_3420 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3289_3289_delayed_14_0_3434 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3297_3297_delayed_14_0_3448 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3305_3305_delayed_14_0_3462 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3313_3313_delayed_14_0_3476 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3321_3321_delayed_14_0_3490 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3329_3329_delayed_14_0_3504 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3337_3337_delayed_14_0_3518 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3345_3345_delayed_14_0_3532 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3353_3353_delayed_14_0_3546 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3361_3361_delayed_14_0_3560 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3369_3369_delayed_14_0_3574 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3377_3377_delayed_14_0_3588 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3385_3385_delayed_14_0_3602 : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_3282_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_3292_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_3158_wire : std_logic_vector(15 downto 0);
    signal MUX_3222_wire : std_logic_vector(15 downto 0);
    signal MUX_3260_wire : std_logic_vector(31 downto 0);
    signal MUX_3274_wire : std_logic_vector(31 downto 0);
    signal NOT_u1_u1_3664_wire : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_3082_3082_delayed_1_0_3198 : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_3430_3430_delayed_1_0_3658 : std_logic_vector(15 downto 0);
    signal UGE_u16_u1_3203_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_3662_wire : std_logic_vector(0 downto 0);
    signal address1_3163 : std_logic_vector(31 downto 0);
    signal address2_3168 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3284_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3284_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3284_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3284_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3284_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3284_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3294_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3294_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3294_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3294_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3294_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3294_root_address : std_logic_vector(13 downto 0);
    signal cb_3151 : std_logic_vector(15 downto 0);
    signal chl_3173 : std_logic_vector(15 downto 0);
    signal chl_change_3205 : std_logic_vector(0 downto 0);
    signal chl_out_3154 : std_logic_vector(15 downto 0);
    signal col_3178 : std_logic_vector(15 downto 0);
    signal continue_flag_3666 : std_logic_vector(0 downto 0);
    signal fetch_addr1_3286 : std_logic_vector(31 downto 0);
    signal fetch_addr1_3390_delayed_8_0_3614 : std_logic_vector(31 downto 0);
    signal fetch_addr2_3296 : std_logic_vector(31 downto 0);
    signal fetch_addr2_3408_delayed_8_0_3635 : std_logic_vector(31 downto 0);
    signal fetch_val1_3300 : std_logic_vector(63 downto 0);
    signal fetch_val2_3304 : std_logic_vector(63 downto 0);
    signal konst_3196_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3208_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3210_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3216_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3219_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3228_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3281_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3291_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3390_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3404_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3418_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3432_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3446_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3460_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3474_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3488_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3502_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3516_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3530_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3544_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3558_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3572_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3586_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3600_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3656_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3670_wire_constant : std_logic_vector(7 downto 0);
    signal location1_3383 : std_logic_vector(2 downto 0);
    signal location2_3387 : std_logic_vector(2 downto 0);
    signal n_address1_3262 : std_logic_vector(31 downto 0);
    signal n_address1_3262_3167_buffered : std_logic_vector(31 downto 0);
    signal n_address2_3276 : std_logic_vector(31 downto 0);
    signal n_address2_3276_3172_buffered : std_logic_vector(31 downto 0);
    signal n_chl_3232 : std_logic_vector(15 downto 0);
    signal n_chl_3232_3177_buffered : std_logic_vector(15 downto 0);
    signal n_col_3213 : std_logic_vector(15 downto 0);
    signal n_col_3213_3182_buffered : std_logic_vector(15 downto 0);
    signal n_row_3224 : std_logic_vector(15 downto 0);
    signal n_row_3224_3187_buffered : std_logic_vector(15 downto 0);
    signal output_data1_3266_delayed_13_0_3395 : std_logic_vector(7 downto 0);
    signal output_data1_3274_delayed_13_0_3409 : std_logic_vector(7 downto 0);
    signal output_data1_3282_delayed_13_0_3423 : std_logic_vector(7 downto 0);
    signal output_data1_3290_delayed_13_0_3437 : std_logic_vector(7 downto 0);
    signal output_data1_3298_delayed_13_0_3451 : std_logic_vector(7 downto 0);
    signal output_data1_3306_delayed_13_0_3465 : std_logic_vector(7 downto 0);
    signal output_data1_3311 : std_logic_vector(7 downto 0);
    signal output_data1_3314_delayed_13_0_3479 : std_logic_vector(7 downto 0);
    signal output_data1_3322_delayed_13_0_3493 : std_logic_vector(7 downto 0);
    signal output_data2_3315 : std_logic_vector(7 downto 0);
    signal output_data2_3330_delayed_13_0_3507 : std_logic_vector(7 downto 0);
    signal output_data2_3338_delayed_13_0_3521 : std_logic_vector(7 downto 0);
    signal output_data2_3346_delayed_13_0_3535 : std_logic_vector(7 downto 0);
    signal output_data2_3354_delayed_13_0_3549 : std_logic_vector(7 downto 0);
    signal output_data2_3362_delayed_13_0_3563 : std_logic_vector(7 downto 0);
    signal output_data2_3370_delayed_13_0_3577 : std_logic_vector(7 downto 0);
    signal output_data2_3378_delayed_13_0_3591 : std_logic_vector(7 downto 0);
    signal output_data2_3386_delayed_13_0_3605 : std_logic_vector(7 downto 0);
    signal output_data_read_3307 : std_logic_vector(15 downto 0);
    signal ptr_deref_3299_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3299_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3299_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3299_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3299_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3303_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3303_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3303_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3303_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3303_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3616_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3616_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3616_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3616_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3616_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3616_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3637_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3637_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3637_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3637_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3637_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3637_word_offset_0 : std_logic_vector(13 downto 0);
    signal rb_3148 : std_logic_vector(15 downto 0);
    signal row_3183 : std_logic_vector(15 downto 0);
    signal row_change_3193 : std_logic_vector(0 downto 0);
    signal row_size_3160 : std_logic_vector(31 downto 0);
    signal tmp1_3241 : std_logic_vector(31 downto 0);
    signal tmp2_3250 : std_logic_vector(31 downto 0);
    signal type_cast_3116_3116_delayed_1_0_3236 : std_logic_vector(31 downto 0);
    signal type_cast_3122_3122_delayed_1_0_3245 : std_logic_vector(31 downto 0);
    signal type_cast_3166_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3171_wire : std_logic_vector(31 downto 0);
    signal type_cast_3176_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3181_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3186_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3254_wire : std_logic_vector(31 downto 0);
    signal type_cast_3266_wire : std_logic_vector(31 downto 0);
    signal type_cast_3283_resized : std_logic_vector(13 downto 0);
    signal type_cast_3283_scaled : std_logic_vector(13 downto 0);
    signal type_cast_3283_wire : std_logic_vector(63 downto 0);
    signal type_cast_3293_resized : std_logic_vector(13 downto 0);
    signal type_cast_3293_scaled : std_logic_vector(13 downto 0);
    signal type_cast_3293_wire : std_logic_vector(63 downto 0);
    signal w11_3319 : std_logic_vector(7 downto 0);
    signal w12_3323 : std_logic_vector(7 downto 0);
    signal w13_3327 : std_logic_vector(7 downto 0);
    signal w14_3331 : std_logic_vector(7 downto 0);
    signal w15_3335 : std_logic_vector(7 downto 0);
    signal w16_3339 : std_logic_vector(7 downto 0);
    signal w17_3343 : std_logic_vector(7 downto 0);
    signal w18_3347 : std_logic_vector(7 downto 0);
    signal w21_3351 : std_logic_vector(7 downto 0);
    signal w22_3355 : std_logic_vector(7 downto 0);
    signal w23_3359 : std_logic_vector(7 downto 0);
    signal w24_3363 : std_logic_vector(7 downto 0);
    signal w25_3367 : std_logic_vector(7 downto 0);
    signal w26_3371 : std_logic_vector(7 downto 0);
    signal w27_3375 : std_logic_vector(7 downto 0);
    signal w28_3379 : std_logic_vector(7 downto 0);
    signal wb11_3401 : std_logic_vector(7 downto 0);
    signal wb12_3415 : std_logic_vector(7 downto 0);
    signal wb13_3429 : std_logic_vector(7 downto 0);
    signal wb14_3443 : std_logic_vector(7 downto 0);
    signal wb15_3457 : std_logic_vector(7 downto 0);
    signal wb16_3471 : std_logic_vector(7 downto 0);
    signal wb17_3485 : std_logic_vector(7 downto 0);
    signal wb18_3499 : std_logic_vector(7 downto 0);
    signal wb21_3513 : std_logic_vector(7 downto 0);
    signal wb22_3527 : std_logic_vector(7 downto 0);
    signal wb23_3541 : std_logic_vector(7 downto 0);
    signal wb24_3555 : std_logic_vector(7 downto 0);
    signal wb25_3569 : std_logic_vector(7 downto 0);
    signal wb26_3583 : std_logic_vector(7 downto 0);
    signal wb27_3597 : std_logic_vector(7 downto 0);
    signal wb28_3611 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_3284_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3284_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3284_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3284_resized_base_address <= "00000000000000";
    array_obj_ref_3294_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3294_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3294_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3294_resized_base_address <= "00000000000000";
    konst_3196_wire_constant <= "0000000000000001";
    konst_3208_wire_constant <= "0000000000000001";
    konst_3210_wire_constant <= "0000000000000001";
    konst_3216_wire_constant <= "0000000000000001";
    konst_3219_wire_constant <= "0000000000000010";
    konst_3228_wire_constant <= "0000000000000001";
    konst_3281_wire_constant <= "00000000000000000000000000000011";
    konst_3291_wire_constant <= "00000000000000000000000000000011";
    konst_3390_wire_constant <= "000";
    konst_3404_wire_constant <= "001";
    konst_3418_wire_constant <= "010";
    konst_3432_wire_constant <= "011";
    konst_3446_wire_constant <= "100";
    konst_3460_wire_constant <= "101";
    konst_3474_wire_constant <= "110";
    konst_3488_wire_constant <= "111";
    konst_3502_wire_constant <= "000";
    konst_3516_wire_constant <= "001";
    konst_3530_wire_constant <= "010";
    konst_3544_wire_constant <= "011";
    konst_3558_wire_constant <= "100";
    konst_3572_wire_constant <= "101";
    konst_3586_wire_constant <= "110";
    konst_3600_wire_constant <= "111";
    konst_3656_wire_constant <= "0000000000000001";
    konst_3670_wire_constant <= "00000001";
    ptr_deref_3299_word_offset_0 <= "00000000000000";
    ptr_deref_3303_word_offset_0 <= "00000000000000";
    ptr_deref_3616_word_offset_0 <= "00000000000000";
    ptr_deref_3637_word_offset_0 <= "00000000000000";
    type_cast_3166_wire_constant <= "00000000000000000000000000000000";
    type_cast_3176_wire_constant <= "0000000000000000";
    type_cast_3181_wire_constant <= "0000000000000001";
    type_cast_3186_wire_constant <= "0000000000000001";
    phi_stmt_3163: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3166_wire_constant & n_address1_3262_3167_buffered;
      req <= phi_stmt_3163_req_0 & phi_stmt_3163_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3163",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3163_ack_0,
          idata => idata,
          odata => address1_3163,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3163
    phi_stmt_3168: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3171_wire & n_address2_3276_3172_buffered;
      req <= phi_stmt_3168_req_0 & phi_stmt_3168_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3168",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3168_ack_0,
          idata => idata,
          odata => address2_3168,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3168
    phi_stmt_3173: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3176_wire_constant & n_chl_3232_3177_buffered;
      req <= phi_stmt_3173_req_0 & phi_stmt_3173_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3173",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3173_ack_0,
          idata => idata,
          odata => chl_3173,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3173
    phi_stmt_3178: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3181_wire_constant & n_col_3213_3182_buffered;
      req <= phi_stmt_3178_req_0 & phi_stmt_3178_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3178",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3178_ack_0,
          idata => idata,
          odata => col_3178,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3178
    phi_stmt_3183: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3186_wire_constant & n_row_3224_3187_buffered;
      req <= phi_stmt_3183_req_0 & phi_stmt_3183_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3183",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3183_ack_0,
          idata => idata,
          odata => row_3183,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3183
    -- flow-through select operator MUX_3212_inst
    n_col_3213 <= konst_3208_wire_constant when (row_change_3193(0) /=  '0') else ADD_u16_u16_3211_wire;
    -- flow-through select operator MUX_3222_inst
    MUX_3222_wire <= ADD_u16_u16_3220_wire when (row_change_3193(0) /=  '0') else row_3183;
    -- flow-through select operator MUX_3223_inst
    n_row_3224 <= konst_3216_wire_constant when (chl_change_3205(0) /=  '0') else MUX_3222_wire;
    -- flow-through select operator MUX_3231_inst
    n_chl_3232 <= ADD_u16_u16_3229_wire when (chl_change_3205(0) /=  '0') else chl_3173;
    -- flow-through select operator MUX_3260_inst
    MUX_3260_wire <= ADD_u32_u32_3258_wire when (row_change_3193(0) /=  '0') else tmp1_3241;
    -- flow-through select operator MUX_3261_inst
    n_address1_3262 <= type_cast_3254_wire when (chl_change_3205(0) /=  '0') else MUX_3260_wire;
    -- flow-through select operator MUX_3274_inst
    MUX_3274_wire <= ADD_u32_u32_3272_wire when (row_change_3193(0) /=  '0') else tmp2_3250;
    -- flow-through select operator MUX_3275_inst
    n_address2_3276 <= ADD_u32_u32_3268_wire when (chl_change_3205(0) /=  '0') else MUX_3274_wire;
    -- flow-through select operator MUX_3400_inst
    wb11_3401 <= output_data1_3266_delayed_13_0_3395 when (EQ_u3_u1_3265_3265_delayed_14_0_3392(0) /=  '0') else w11_3319;
    -- flow-through select operator MUX_3414_inst
    wb12_3415 <= output_data1_3274_delayed_13_0_3409 when (EQ_u3_u1_3273_3273_delayed_14_0_3406(0) /=  '0') else w12_3323;
    -- flow-through select operator MUX_3428_inst
    wb13_3429 <= output_data1_3282_delayed_13_0_3423 when (EQ_u3_u1_3281_3281_delayed_14_0_3420(0) /=  '0') else w13_3327;
    -- flow-through select operator MUX_3442_inst
    wb14_3443 <= output_data1_3290_delayed_13_0_3437 when (EQ_u3_u1_3289_3289_delayed_14_0_3434(0) /=  '0') else w14_3331;
    -- flow-through select operator MUX_3456_inst
    wb15_3457 <= output_data1_3298_delayed_13_0_3451 when (EQ_u3_u1_3297_3297_delayed_14_0_3448(0) /=  '0') else w15_3335;
    -- flow-through select operator MUX_3470_inst
    wb16_3471 <= output_data1_3306_delayed_13_0_3465 when (EQ_u3_u1_3305_3305_delayed_14_0_3462(0) /=  '0') else w16_3339;
    -- flow-through select operator MUX_3484_inst
    wb17_3485 <= output_data1_3314_delayed_13_0_3479 when (EQ_u3_u1_3313_3313_delayed_14_0_3476(0) /=  '0') else w17_3343;
    -- flow-through select operator MUX_3498_inst
    wb18_3499 <= output_data1_3322_delayed_13_0_3493 when (EQ_u3_u1_3321_3321_delayed_14_0_3490(0) /=  '0') else w18_3347;
    -- flow-through select operator MUX_3512_inst
    wb21_3513 <= output_data2_3330_delayed_13_0_3507 when (EQ_u3_u1_3329_3329_delayed_14_0_3504(0) /=  '0') else w21_3351;
    -- flow-through select operator MUX_3526_inst
    wb22_3527 <= output_data2_3338_delayed_13_0_3521 when (EQ_u3_u1_3337_3337_delayed_14_0_3518(0) /=  '0') else w22_3355;
    -- flow-through select operator MUX_3540_inst
    wb23_3541 <= output_data2_3346_delayed_13_0_3535 when (EQ_u3_u1_3345_3345_delayed_14_0_3532(0) /=  '0') else w23_3359;
    -- flow-through select operator MUX_3554_inst
    wb24_3555 <= output_data2_3354_delayed_13_0_3549 when (EQ_u3_u1_3353_3353_delayed_14_0_3546(0) /=  '0') else w24_3363;
    -- flow-through select operator MUX_3568_inst
    wb25_3569 <= output_data2_3362_delayed_13_0_3563 when (EQ_u3_u1_3361_3361_delayed_14_0_3560(0) /=  '0') else w25_3367;
    -- flow-through select operator MUX_3582_inst
    wb26_3583 <= output_data2_3370_delayed_13_0_3577 when (EQ_u3_u1_3369_3369_delayed_14_0_3574(0) /=  '0') else w26_3371;
    -- flow-through select operator MUX_3596_inst
    wb27_3597 <= output_data2_3378_delayed_13_0_3591 when (EQ_u3_u1_3377_3377_delayed_14_0_3588(0) /=  '0') else w27_3375;
    -- flow-through select operator MUX_3610_inst
    wb28_3611 <= output_data2_3386_delayed_13_0_3605 when (EQ_u3_u1_3385_3385_delayed_14_0_3602(0) /=  '0') else w28_3379;
    slice_3310_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3310_inst_req_0;
      slice_3310_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3310_inst_req_1;
      slice_3310_inst_ack_1<= update_ack(0);
      slice_3310_inst: SliceSplitProtocol generic map(name => "slice_3310_inst", in_data_width => 16, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => output_data_read_3307, dout => output_data1_3311, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3314_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3314_inst_req_0;
      slice_3314_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3314_inst_req_1;
      slice_3314_inst_ack_1<= update_ack(0);
      slice_3314_inst: SliceSplitProtocol generic map(name => "slice_3314_inst", in_data_width => 16, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => output_data_read_3307, dout => output_data2_3315, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3318_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3318_inst_req_0;
      slice_3318_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3318_inst_req_1;
      slice_3318_inst_ack_1<= update_ack(0);
      slice_3318_inst: SliceSplitProtocol generic map(name => "slice_3318_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3300, dout => w11_3319, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3322_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3322_inst_req_0;
      slice_3322_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3322_inst_req_1;
      slice_3322_inst_ack_1<= update_ack(0);
      slice_3322_inst: SliceSplitProtocol generic map(name => "slice_3322_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3300, dout => w12_3323, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3326_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3326_inst_req_0;
      slice_3326_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3326_inst_req_1;
      slice_3326_inst_ack_1<= update_ack(0);
      slice_3326_inst: SliceSplitProtocol generic map(name => "slice_3326_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3300, dout => w13_3327, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3330_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3330_inst_req_0;
      slice_3330_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3330_inst_req_1;
      slice_3330_inst_ack_1<= update_ack(0);
      slice_3330_inst: SliceSplitProtocol generic map(name => "slice_3330_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3300, dout => w14_3331, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3334_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3334_inst_req_0;
      slice_3334_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3334_inst_req_1;
      slice_3334_inst_ack_1<= update_ack(0);
      slice_3334_inst: SliceSplitProtocol generic map(name => "slice_3334_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3300, dout => w15_3335, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3338_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3338_inst_req_0;
      slice_3338_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3338_inst_req_1;
      slice_3338_inst_ack_1<= update_ack(0);
      slice_3338_inst: SliceSplitProtocol generic map(name => "slice_3338_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3300, dout => w16_3339, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3342_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3342_inst_req_0;
      slice_3342_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3342_inst_req_1;
      slice_3342_inst_ack_1<= update_ack(0);
      slice_3342_inst: SliceSplitProtocol generic map(name => "slice_3342_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3300, dout => w17_3343, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3346_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3346_inst_req_0;
      slice_3346_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3346_inst_req_1;
      slice_3346_inst_ack_1<= update_ack(0);
      slice_3346_inst: SliceSplitProtocol generic map(name => "slice_3346_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3300, dout => w18_3347, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3350_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3350_inst_req_0;
      slice_3350_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3350_inst_req_1;
      slice_3350_inst_ack_1<= update_ack(0);
      slice_3350_inst: SliceSplitProtocol generic map(name => "slice_3350_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3304, dout => w21_3351, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3354_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3354_inst_req_0;
      slice_3354_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3354_inst_req_1;
      slice_3354_inst_ack_1<= update_ack(0);
      slice_3354_inst: SliceSplitProtocol generic map(name => "slice_3354_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3304, dout => w22_3355, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3358_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3358_inst_req_0;
      slice_3358_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3358_inst_req_1;
      slice_3358_inst_ack_1<= update_ack(0);
      slice_3358_inst: SliceSplitProtocol generic map(name => "slice_3358_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3304, dout => w23_3359, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3362_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3362_inst_req_0;
      slice_3362_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3362_inst_req_1;
      slice_3362_inst_ack_1<= update_ack(0);
      slice_3362_inst: SliceSplitProtocol generic map(name => "slice_3362_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3304, dout => w24_3363, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3366_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3366_inst_req_0;
      slice_3366_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3366_inst_req_1;
      slice_3366_inst_ack_1<= update_ack(0);
      slice_3366_inst: SliceSplitProtocol generic map(name => "slice_3366_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3304, dout => w25_3367, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3370_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3370_inst_req_0;
      slice_3370_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3370_inst_req_1;
      slice_3370_inst_ack_1<= update_ack(0);
      slice_3370_inst: SliceSplitProtocol generic map(name => "slice_3370_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3304, dout => w26_3371, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3374_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3374_inst_req_0;
      slice_3374_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3374_inst_req_1;
      slice_3374_inst_ack_1<= update_ack(0);
      slice_3374_inst: SliceSplitProtocol generic map(name => "slice_3374_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3304, dout => w27_3375, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3378_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3378_inst_req_0;
      slice_3378_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3378_inst_req_1;
      slice_3378_inst_ack_1<= update_ack(0);
      slice_3378_inst: SliceSplitProtocol generic map(name => "slice_3378_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3304, dout => w28_3379, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_fetch_addr1_3390_delayed_8_0_3612_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_addr1_3390_delayed_8_0_3612_inst_req_0;
      W_fetch_addr1_3390_delayed_8_0_3612_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_addr1_3390_delayed_8_0_3612_inst_req_1;
      W_fetch_addr1_3390_delayed_8_0_3612_inst_ack_1<= rack(0);
      W_fetch_addr1_3390_delayed_8_0_3612_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_addr1_3390_delayed_8_0_3612_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_addr1_3286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_3390_delayed_8_0_3614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_addr2_3408_delayed_8_0_3633_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_addr2_3408_delayed_8_0_3633_inst_req_0;
      W_fetch_addr2_3408_delayed_8_0_3633_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_addr2_3408_delayed_8_0_3633_inst_req_1;
      W_fetch_addr2_3408_delayed_8_0_3633_inst_ack_1<= rack(0);
      W_fetch_addr2_3408_delayed_8_0_3633_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_addr2_3408_delayed_8_0_3633_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_addr2_3296,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_3408_delayed_8_0_3635,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3266_delayed_13_0_3393_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3266_delayed_13_0_3393_inst_req_0;
      W_output_data1_3266_delayed_13_0_3393_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3266_delayed_13_0_3393_inst_req_1;
      W_output_data1_3266_delayed_13_0_3393_inst_ack_1<= rack(0);
      W_output_data1_3266_delayed_13_0_3393_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3266_delayed_13_0_3393_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3266_delayed_13_0_3395,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3274_delayed_13_0_3407_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3274_delayed_13_0_3407_inst_req_0;
      W_output_data1_3274_delayed_13_0_3407_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3274_delayed_13_0_3407_inst_req_1;
      W_output_data1_3274_delayed_13_0_3407_inst_ack_1<= rack(0);
      W_output_data1_3274_delayed_13_0_3407_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3274_delayed_13_0_3407_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3274_delayed_13_0_3409,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3282_delayed_13_0_3421_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3282_delayed_13_0_3421_inst_req_0;
      W_output_data1_3282_delayed_13_0_3421_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3282_delayed_13_0_3421_inst_req_1;
      W_output_data1_3282_delayed_13_0_3421_inst_ack_1<= rack(0);
      W_output_data1_3282_delayed_13_0_3421_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3282_delayed_13_0_3421_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3282_delayed_13_0_3423,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3290_delayed_13_0_3435_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3290_delayed_13_0_3435_inst_req_0;
      W_output_data1_3290_delayed_13_0_3435_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3290_delayed_13_0_3435_inst_req_1;
      W_output_data1_3290_delayed_13_0_3435_inst_ack_1<= rack(0);
      W_output_data1_3290_delayed_13_0_3435_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3290_delayed_13_0_3435_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3290_delayed_13_0_3437,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3298_delayed_13_0_3449_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3298_delayed_13_0_3449_inst_req_0;
      W_output_data1_3298_delayed_13_0_3449_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3298_delayed_13_0_3449_inst_req_1;
      W_output_data1_3298_delayed_13_0_3449_inst_ack_1<= rack(0);
      W_output_data1_3298_delayed_13_0_3449_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3298_delayed_13_0_3449_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3298_delayed_13_0_3451,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3306_delayed_13_0_3463_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3306_delayed_13_0_3463_inst_req_0;
      W_output_data1_3306_delayed_13_0_3463_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3306_delayed_13_0_3463_inst_req_1;
      W_output_data1_3306_delayed_13_0_3463_inst_ack_1<= rack(0);
      W_output_data1_3306_delayed_13_0_3463_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3306_delayed_13_0_3463_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3306_delayed_13_0_3465,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3314_delayed_13_0_3477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3314_delayed_13_0_3477_inst_req_0;
      W_output_data1_3314_delayed_13_0_3477_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3314_delayed_13_0_3477_inst_req_1;
      W_output_data1_3314_delayed_13_0_3477_inst_ack_1<= rack(0);
      W_output_data1_3314_delayed_13_0_3477_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3314_delayed_13_0_3477_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3314_delayed_13_0_3479,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3322_delayed_13_0_3491_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3322_delayed_13_0_3491_inst_req_0;
      W_output_data1_3322_delayed_13_0_3491_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3322_delayed_13_0_3491_inst_req_1;
      W_output_data1_3322_delayed_13_0_3491_inst_ack_1<= rack(0);
      W_output_data1_3322_delayed_13_0_3491_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3322_delayed_13_0_3491_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3311,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3322_delayed_13_0_3493,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3330_delayed_13_0_3505_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3330_delayed_13_0_3505_inst_req_0;
      W_output_data2_3330_delayed_13_0_3505_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3330_delayed_13_0_3505_inst_req_1;
      W_output_data2_3330_delayed_13_0_3505_inst_ack_1<= rack(0);
      W_output_data2_3330_delayed_13_0_3505_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3330_delayed_13_0_3505_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3330_delayed_13_0_3507,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3338_delayed_13_0_3519_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3338_delayed_13_0_3519_inst_req_0;
      W_output_data2_3338_delayed_13_0_3519_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3338_delayed_13_0_3519_inst_req_1;
      W_output_data2_3338_delayed_13_0_3519_inst_ack_1<= rack(0);
      W_output_data2_3338_delayed_13_0_3519_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3338_delayed_13_0_3519_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3338_delayed_13_0_3521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3346_delayed_13_0_3533_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3346_delayed_13_0_3533_inst_req_0;
      W_output_data2_3346_delayed_13_0_3533_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3346_delayed_13_0_3533_inst_req_1;
      W_output_data2_3346_delayed_13_0_3533_inst_ack_1<= rack(0);
      W_output_data2_3346_delayed_13_0_3533_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3346_delayed_13_0_3533_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3346_delayed_13_0_3535,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3354_delayed_13_0_3547_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3354_delayed_13_0_3547_inst_req_0;
      W_output_data2_3354_delayed_13_0_3547_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3354_delayed_13_0_3547_inst_req_1;
      W_output_data2_3354_delayed_13_0_3547_inst_ack_1<= rack(0);
      W_output_data2_3354_delayed_13_0_3547_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3354_delayed_13_0_3547_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3354_delayed_13_0_3549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3362_delayed_13_0_3561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3362_delayed_13_0_3561_inst_req_0;
      W_output_data2_3362_delayed_13_0_3561_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3362_delayed_13_0_3561_inst_req_1;
      W_output_data2_3362_delayed_13_0_3561_inst_ack_1<= rack(0);
      W_output_data2_3362_delayed_13_0_3561_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3362_delayed_13_0_3561_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3362_delayed_13_0_3563,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3370_delayed_13_0_3575_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3370_delayed_13_0_3575_inst_req_0;
      W_output_data2_3370_delayed_13_0_3575_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3370_delayed_13_0_3575_inst_req_1;
      W_output_data2_3370_delayed_13_0_3575_inst_ack_1<= rack(0);
      W_output_data2_3370_delayed_13_0_3575_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3370_delayed_13_0_3575_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3370_delayed_13_0_3577,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3378_delayed_13_0_3589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3378_delayed_13_0_3589_inst_req_0;
      W_output_data2_3378_delayed_13_0_3589_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3378_delayed_13_0_3589_inst_req_1;
      W_output_data2_3378_delayed_13_0_3589_inst_ack_1<= rack(0);
      W_output_data2_3378_delayed_13_0_3589_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3378_delayed_13_0_3589_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3378_delayed_13_0_3591,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3386_delayed_13_0_3603_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3386_delayed_13_0_3603_inst_req_0;
      W_output_data2_3386_delayed_13_0_3603_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3386_delayed_13_0_3603_inst_req_1;
      W_output_data2_3386_delayed_13_0_3603_inst_ack_1<= rack(0);
      W_output_data2_3386_delayed_13_0_3603_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3386_delayed_13_0_3603_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3386_delayed_13_0_3605,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3285_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3285_final_reg_req_0;
      addr_of_3285_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3285_final_reg_req_1;
      addr_of_3285_final_reg_ack_1<= rack(0);
      addr_of_3285_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3285_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3284_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_3286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3295_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3295_final_reg_req_0;
      addr_of_3295_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3295_final_reg_req_1;
      addr_of_3295_final_reg_ack_1<= rack(0);
      addr_of_3295_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3295_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3294_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_3296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address1_3262_3167_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address1_3262_3167_buf_req_0;
      n_address1_3262_3167_buf_ack_0<= wack(0);
      rreq(0) <= n_address1_3262_3167_buf_req_1;
      n_address1_3262_3167_buf_ack_1<= rack(0);
      n_address1_3262_3167_buf : InterlockBuffer generic map ( -- 
        name => "n_address1_3262_3167_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address1_3262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address1_3262_3167_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address2_3276_3172_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address2_3276_3172_buf_req_0;
      n_address2_3276_3172_buf_ack_0<= wack(0);
      rreq(0) <= n_address2_3276_3172_buf_req_1;
      n_address2_3276_3172_buf_ack_1<= rack(0);
      n_address2_3276_3172_buf : InterlockBuffer generic map ( -- 
        name => "n_address2_3276_3172_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address2_3276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address2_3276_3172_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_3232_3177_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_3232_3177_buf_req_0;
      n_chl_3232_3177_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_3232_3177_buf_req_1;
      n_chl_3232_3177_buf_ack_1<= rack(0);
      n_chl_3232_3177_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_3232_3177_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_3232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_3232_3177_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_3213_3182_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_3213_3182_buf_req_0;
      n_col_3213_3182_buf_ack_0<= wack(0);
      rreq(0) <= n_col_3213_3182_buf_req_1;
      n_col_3213_3182_buf_ack_1<= rack(0);
      n_col_3213_3182_buf : InterlockBuffer generic map ( -- 
        name => "n_col_3213_3182_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_3213,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_3213_3182_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_3224_3187_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_3224_3187_buf_req_0;
      n_row_3224_3187_buf_ack_0<= wack(0);
      rreq(0) <= n_row_3224_3187_buf_req_1;
      n_row_3224_3187_buf_ack_1<= rack(0);
      n_row_3224_3187_buf : InterlockBuffer generic map ( -- 
        name => "n_row_3224_3187_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_3224,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_3224_3187_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3159_inst
    process(MUL_u16_u16_3158_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_3158_wire(15 downto 0);
      row_size_3160 <= tmp_var; -- 
    end process;
    type_cast_3171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3171_inst_req_0;
      type_cast_3171_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3171_inst_req_1;
      type_cast_3171_inst_ack_1<= rack(0);
      type_cast_3171_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3171_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => row_size_3160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3171_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3235_inst_req_0;
      type_cast_3235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3235_inst_req_1;
      type_cast_3235_inst_ack_1<= rack(0);
      type_cast_3235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3235_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chl_out_3154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3116_3116_delayed_1_0_3236,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3244_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3244_inst_req_0;
      type_cast_3244_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3244_inst_req_1;
      type_cast_3244_inst_ack_1<= rack(0);
      type_cast_3244_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3244_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chl_out_3154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3122_3122_delayed_1_0_3245,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3254_inst
    process(n_chl_3232) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_chl_3232(15 downto 0);
      type_cast_3254_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3266_inst
    process(n_chl_3232) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_chl_3232(15 downto 0);
      type_cast_3266_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3283_inst
    process(LSHR_u32_u32_3282_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_3282_wire(31 downto 0);
      type_cast_3283_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3293_inst
    process(LSHR_u32_u32_3292_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_3292_wire(31 downto 0);
      type_cast_3293_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3382_inst
    process(address1_3163) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 2 downto 0) := address1_3163(2 downto 0);
      location1_3383 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3386_inst
    process(address2_3168) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 2 downto 0) := address2_3168(2 downto 0);
      location2_3387 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_3284_index_1_rename
    process(type_cast_3283_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3283_resized;
      ov(13 downto 0) := iv;
      type_cast_3283_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3284_index_1_resize
    process(type_cast_3283_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3283_wire;
      ov := iv(13 downto 0);
      type_cast_3283_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3284_root_address_inst
    process(array_obj_ref_3284_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3284_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3284_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3294_index_1_rename
    process(type_cast_3293_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3293_resized;
      ov(13 downto 0) := iv;
      type_cast_3293_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3294_index_1_resize
    process(type_cast_3293_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3293_wire;
      ov := iv(13 downto 0);
      type_cast_3293_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3294_root_address_inst
    process(array_obj_ref_3294_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3294_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3294_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3299_addr_0
    process(ptr_deref_3299_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3299_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3299_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3299_base_resize
    process(fetch_addr1_3286) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_3286;
      ov := iv(13 downto 0);
      ptr_deref_3299_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3299_gather_scatter
    process(ptr_deref_3299_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3299_data_0;
      ov(63 downto 0) := iv;
      fetch_val1_3300 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3299_root_address_inst
    process(ptr_deref_3299_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3299_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3299_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3303_addr_0
    process(ptr_deref_3303_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3303_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3303_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3303_base_resize
    process(fetch_addr2_3296) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_3296;
      ov := iv(13 downto 0);
      ptr_deref_3303_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3303_gather_scatter
    process(ptr_deref_3303_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3303_data_0;
      ov(63 downto 0) := iv;
      fetch_val2_3304 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3303_root_address_inst
    process(ptr_deref_3303_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3303_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3303_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3616_addr_0
    process(ptr_deref_3616_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3616_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3616_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3616_base_resize
    process(fetch_addr1_3390_delayed_8_0_3614) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_3390_delayed_8_0_3614;
      ov := iv(13 downto 0);
      ptr_deref_3616_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3616_gather_scatter
    process(CONCAT_u32_u64_3631_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_3631_wire;
      ov(63 downto 0) := iv;
      ptr_deref_3616_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3616_root_address_inst
    process(ptr_deref_3616_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3616_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3616_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3637_addr_0
    process(ptr_deref_3637_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3637_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3637_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3637_base_resize
    process(fetch_addr2_3408_delayed_8_0_3635) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_3408_delayed_8_0_3635;
      ov := iv(13 downto 0);
      ptr_deref_3637_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3637_gather_scatter
    process(CONCAT_u32_u64_3652_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_3652_wire;
      ov(63 downto 0) := iv;
      ptr_deref_3637_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3637_root_address_inst
    process(ptr_deref_3637_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3637_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3637_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_3161_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_3666;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_3161_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_3161_branch_req_0,
          ack0 => do_while_stmt_3161_branch_ack_0,
          ack1 => do_while_stmt_3161_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3211_inst
    process(col_3178) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_3178, konst_3210_wire_constant, tmp_var);
      ADD_u16_u16_3211_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3220_inst
    process(row_3183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_3183, konst_3219_wire_constant, tmp_var);
      ADD_u16_u16_3220_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3229_inst
    process(chl_3173) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_3173, konst_3228_wire_constant, tmp_var);
      ADD_u16_u16_3229_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3240_inst
    process(address1_3163, type_cast_3116_3116_delayed_1_0_3236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address1_3163, type_cast_3116_3116_delayed_1_0_3236, tmp_var);
      tmp1_3241 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3249_inst
    process(address2_3168, type_cast_3122_3122_delayed_1_0_3245) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address2_3168, type_cast_3122_3122_delayed_1_0_3245, tmp_var);
      tmp2_3250 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3258_inst
    process(tmp1_3241, row_size_3160) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_3241, row_size_3160, tmp_var);
      ADD_u32_u32_3258_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3268_inst
    process(type_cast_3266_wire, row_size_3160) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_3266_wire, row_size_3160, tmp_var);
      ADD_u32_u32_3268_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3272_inst
    process(tmp2_3250, row_size_3160) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp2_3250, row_size_3160, tmp_var);
      ADD_u32_u32_3272_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3204_inst
    process(row_change_3193, UGE_u16_u1_3203_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(row_change_3193, UGE_u16_u1_3203_wire, tmp_var);
      chl_change_3205 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3623_inst
    process(CONCAT_u8_u16_3619_wire, CONCAT_u8_u16_3622_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_3619_wire, CONCAT_u8_u16_3622_wire, tmp_var);
      CONCAT_u16_u32_3623_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3630_inst
    process(CONCAT_u8_u16_3626_wire, CONCAT_u8_u16_3629_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_3626_wire, CONCAT_u8_u16_3629_wire, tmp_var);
      CONCAT_u16_u32_3630_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3644_inst
    process(CONCAT_u8_u16_3640_wire, CONCAT_u8_u16_3643_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_3640_wire, CONCAT_u8_u16_3643_wire, tmp_var);
      CONCAT_u16_u32_3644_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3651_inst
    process(CONCAT_u8_u16_3647_wire, CONCAT_u8_u16_3650_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_3647_wire, CONCAT_u8_u16_3650_wire, tmp_var);
      CONCAT_u16_u32_3651_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : CONCAT_u32_u64_3631_inst 
    ApConcat_group_13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_3623_wire & CONCAT_u16_u32_3630_wire;
      CONCAT_u32_u64_3631_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_3631_inst_req_0;
      CONCAT_u32_u64_3631_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_3631_inst_req_1;
      CONCAT_u32_u64_3631_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_13_gI: SplitGuardInterface generic map(name => "ApConcat_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : CONCAT_u32_u64_3652_inst 
    ApConcat_group_14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_3644_wire & CONCAT_u16_u32_3651_wire;
      CONCAT_u32_u64_3652_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_3652_inst_req_0;
      CONCAT_u32_u64_3652_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_3652_inst_req_1;
      CONCAT_u32_u64_3652_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_14_gI: SplitGuardInterface generic map(name => "ApConcat_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- binary operator CONCAT_u8_u16_3619_inst
    process(wb11_3401, wb12_3415) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb11_3401, wb12_3415, tmp_var);
      CONCAT_u8_u16_3619_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3622_inst
    process(wb13_3429, wb14_3443) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb13_3429, wb14_3443, tmp_var);
      CONCAT_u8_u16_3622_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3626_inst
    process(wb15_3457, wb16_3471) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb15_3457, wb16_3471, tmp_var);
      CONCAT_u8_u16_3626_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3629_inst
    process(wb17_3485, wb18_3499) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb17_3485, wb18_3499, tmp_var);
      CONCAT_u8_u16_3629_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3640_inst
    process(wb21_3513, wb22_3527) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb21_3513, wb22_3527, tmp_var);
      CONCAT_u8_u16_3640_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3643_inst
    process(wb23_3541, wb24_3555) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb23_3541, wb24_3555, tmp_var);
      CONCAT_u8_u16_3643_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3647_inst
    process(wb25_3569, wb26_3583) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb25_3569, wb26_3583, tmp_var);
      CONCAT_u8_u16_3647_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3650_inst
    process(wb27_3597, wb28_3611) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb27_3597, wb28_3611, tmp_var);
      CONCAT_u8_u16_3650_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_3192_inst
    process(col_3178, cb_3151) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_3178, cb_3151, tmp_var);
      row_change_3193 <= tmp_var; --
    end process;
    -- shared split operator group (24) : EQ_u3_u1_3391_inst 
    ApIntEq_group_24: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3383;
      EQ_u3_u1_3265_3265_delayed_14_0_3392 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3391_inst_req_0;
      EQ_u3_u1_3391_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3391_inst_req_1;
      EQ_u3_u1_3391_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_24_gI: SplitGuardInterface generic map(name => "ApIntEq_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : EQ_u3_u1_3405_inst 
    ApIntEq_group_25: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3383;
      EQ_u3_u1_3273_3273_delayed_14_0_3406 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3405_inst_req_0;
      EQ_u3_u1_3405_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3405_inst_req_1;
      EQ_u3_u1_3405_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_25_gI: SplitGuardInterface generic map(name => "ApIntEq_group_25_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_25",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "001",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : EQ_u3_u1_3419_inst 
    ApIntEq_group_26: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3383;
      EQ_u3_u1_3281_3281_delayed_14_0_3420 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3419_inst_req_0;
      EQ_u3_u1_3419_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3419_inst_req_1;
      EQ_u3_u1_3419_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_26_gI: SplitGuardInterface generic map(name => "ApIntEq_group_26_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_26",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "010",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : EQ_u3_u1_3433_inst 
    ApIntEq_group_27: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3383;
      EQ_u3_u1_3289_3289_delayed_14_0_3434 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3433_inst_req_0;
      EQ_u3_u1_3433_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3433_inst_req_1;
      EQ_u3_u1_3433_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_27_gI: SplitGuardInterface generic map(name => "ApIntEq_group_27_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "011",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : EQ_u3_u1_3447_inst 
    ApIntEq_group_28: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3383;
      EQ_u3_u1_3297_3297_delayed_14_0_3448 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3447_inst_req_0;
      EQ_u3_u1_3447_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3447_inst_req_1;
      EQ_u3_u1_3447_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_28_gI: SplitGuardInterface generic map(name => "ApIntEq_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "100",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : EQ_u3_u1_3461_inst 
    ApIntEq_group_29: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3383;
      EQ_u3_u1_3305_3305_delayed_14_0_3462 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3461_inst_req_0;
      EQ_u3_u1_3461_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3461_inst_req_1;
      EQ_u3_u1_3461_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_29_gI: SplitGuardInterface generic map(name => "ApIntEq_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "101",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : EQ_u3_u1_3475_inst 
    ApIntEq_group_30: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3383;
      EQ_u3_u1_3313_3313_delayed_14_0_3476 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3475_inst_req_0;
      EQ_u3_u1_3475_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3475_inst_req_1;
      EQ_u3_u1_3475_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_30_gI: SplitGuardInterface generic map(name => "ApIntEq_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "110",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : EQ_u3_u1_3489_inst 
    ApIntEq_group_31: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3383;
      EQ_u3_u1_3321_3321_delayed_14_0_3490 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3489_inst_req_0;
      EQ_u3_u1_3489_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3489_inst_req_1;
      EQ_u3_u1_3489_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_31_gI: SplitGuardInterface generic map(name => "ApIntEq_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "111",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : EQ_u3_u1_3503_inst 
    ApIntEq_group_32: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3387;
      EQ_u3_u1_3329_3329_delayed_14_0_3504 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3503_inst_req_0;
      EQ_u3_u1_3503_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3503_inst_req_1;
      EQ_u3_u1_3503_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_32_gI: SplitGuardInterface generic map(name => "ApIntEq_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : EQ_u3_u1_3517_inst 
    ApIntEq_group_33: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3387;
      EQ_u3_u1_3337_3337_delayed_14_0_3518 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3517_inst_req_0;
      EQ_u3_u1_3517_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3517_inst_req_1;
      EQ_u3_u1_3517_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_33_gI: SplitGuardInterface generic map(name => "ApIntEq_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "001",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : EQ_u3_u1_3531_inst 
    ApIntEq_group_34: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3387;
      EQ_u3_u1_3345_3345_delayed_14_0_3532 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3531_inst_req_0;
      EQ_u3_u1_3531_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3531_inst_req_1;
      EQ_u3_u1_3531_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_34_gI: SplitGuardInterface generic map(name => "ApIntEq_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "010",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : EQ_u3_u1_3545_inst 
    ApIntEq_group_35: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3387;
      EQ_u3_u1_3353_3353_delayed_14_0_3546 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3545_inst_req_0;
      EQ_u3_u1_3545_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3545_inst_req_1;
      EQ_u3_u1_3545_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_35_gI: SplitGuardInterface generic map(name => "ApIntEq_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "011",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : EQ_u3_u1_3559_inst 
    ApIntEq_group_36: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3387;
      EQ_u3_u1_3361_3361_delayed_14_0_3560 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3559_inst_req_0;
      EQ_u3_u1_3559_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3559_inst_req_1;
      EQ_u3_u1_3559_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_36_gI: SplitGuardInterface generic map(name => "ApIntEq_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "100",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : EQ_u3_u1_3573_inst 
    ApIntEq_group_37: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3387;
      EQ_u3_u1_3369_3369_delayed_14_0_3574 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3573_inst_req_0;
      EQ_u3_u1_3573_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3573_inst_req_1;
      EQ_u3_u1_3573_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_37_gI: SplitGuardInterface generic map(name => "ApIntEq_group_37_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "101",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : EQ_u3_u1_3587_inst 
    ApIntEq_group_38: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3387;
      EQ_u3_u1_3377_3377_delayed_14_0_3588 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3587_inst_req_0;
      EQ_u3_u1_3587_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3587_inst_req_1;
      EQ_u3_u1_3587_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_38_gI: SplitGuardInterface generic map(name => "ApIntEq_group_38_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "110",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : EQ_u3_u1_3601_inst 
    ApIntEq_group_39: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3387;
      EQ_u3_u1_3385_3385_delayed_14_0_3602 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3601_inst_req_0;
      EQ_u3_u1_3601_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3601_inst_req_1;
      EQ_u3_u1_3601_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_39_gI: SplitGuardInterface generic map(name => "ApIntEq_group_39_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_39",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "111",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- binary operator LSHR_u32_u32_3282_inst
    process(address1_3163) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address1_3163, konst_3281_wire_constant, tmp_var);
      LSHR_u32_u32_3282_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3292_inst
    process(address2_3168) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address2_3168, konst_3291_wire_constant, tmp_var);
      LSHR_u32_u32_3292_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3158_inst
    process(chl_out_3154, cb_3151) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_out_3154, cb_3151, tmp_var);
      MUL_u16_u16_3158_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_3664_inst
    process(chl_change_3205) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", chl_change_3205, tmp_var);
      NOT_u1_u1_3664_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_3665_inst
    process(ULT_u16_u1_3662_wire, NOT_u1_u1_3664_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ULT_u16_u1_3662_wire, NOT_u1_u1_3664_wire, tmp_var);
      continue_flag_3666 <= tmp_var; --
    end process;
    -- shared split operator group (45) : SUB_u16_u16_3197_inst 
    ApIntSub_group_45: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rb_3148;
      SUB_u16_u16_3082_3082_delayed_1_0_3198 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_3197_inst_req_0;
      SUB_u16_u16_3197_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_3197_inst_req_1;
      SUB_u16_u16_3197_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_45_gI: SplitGuardInterface generic map(name => "ApIntSub_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : SUB_u16_u16_3657_inst 
    ApIntSub_group_46: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= chl_out_3154;
      SUB_u16_u16_3430_3430_delayed_1_0_3658 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_3657_inst_req_0;
      SUB_u16_u16_3657_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_3657_inst_req_1;
      SUB_u16_u16_3657_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_46_gI: SplitGuardInterface generic map(name => "ApIntSub_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- binary operator UGE_u16_u1_3203_inst
    process(row_3183, SUB_u16_u16_3082_3082_delayed_1_0_3198) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(row_3183, SUB_u16_u16_3082_3082_delayed_1_0_3198, tmp_var);
      UGE_u16_u1_3203_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_3662_inst
    process(chl_3173, SUB_u16_u16_3430_3430_delayed_1_0_3658) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(chl_3173, SUB_u16_u16_3430_3430_delayed_1_0_3658, tmp_var);
      ULT_u16_u1_3662_wire <= tmp_var; --
    end process;
    -- shared split operator group (49) : array_obj_ref_3284_index_offset 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3283_scaled;
      array_obj_ref_3284_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3284_index_offset_req_0;
      array_obj_ref_3284_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3284_index_offset_req_1;
      array_obj_ref_3284_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_49_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : array_obj_ref_3294_index_offset 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3293_scaled;
      array_obj_ref_3294_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3294_index_offset_req_0;
      array_obj_ref_3294_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3294_index_offset_req_1;
      array_obj_ref_3294_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared load operator group (0) : ptr_deref_3299_load_0 ptr_deref_3303_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3299_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3303_load_0_req_0;
      ptr_deref_3299_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3303_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3299_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3303_load_0_req_1;
      ptr_deref_3299_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3303_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3299_word_address_0 & ptr_deref_3303_word_address_0;
      ptr_deref_3299_data_0 <= data_out(127 downto 64);
      ptr_deref_3303_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_3616_store_0 ptr_deref_3637_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3616_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3637_store_0_req_0;
      ptr_deref_3616_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3637_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3616_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3637_store_0_req_1;
      ptr_deref_3616_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3637_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3616_word_address_0 & ptr_deref_3637_word_address_0;
      data_in <= ptr_deref_3616_data_0 & ptr_deref_3637_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_output_pipe_3147_inst RPIPE_output_pipe_3150_inst RPIPE_output_pipe_3153_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(47 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 2 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= RPIPE_output_pipe_3147_inst_req_0;
      reqL_unguarded(1) <= RPIPE_output_pipe_3150_inst_req_0;
      reqL_unguarded(0) <= RPIPE_output_pipe_3153_inst_req_0;
      RPIPE_output_pipe_3147_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_output_pipe_3150_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_output_pipe_3153_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= RPIPE_output_pipe_3147_inst_req_1;
      reqR_unguarded(1) <= RPIPE_output_pipe_3150_inst_req_1;
      reqR_unguarded(0) <= RPIPE_output_pipe_3153_inst_req_1;
      RPIPE_output_pipe_3147_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_output_pipe_3150_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_output_pipe_3153_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      rb_3148 <= data_out(47 downto 32);
      cb_3151 <= data_out(31 downto 16);
      chl_out_3154 <= data_out(15 downto 0);
      output_pipe_read_0_gI: SplitGuardInterface generic map(name => "output_pipe_read_0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      output_pipe_read_0: InputPortRevised -- 
        generic map ( name => "output_pipe_read_0", data_width => 16,  num_reqs => 3,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => output_pipe_pipe_read_req(1),
          oack => output_pipe_pipe_read_ack(1),
          odata => output_pipe_pipe_read_data(31 downto 16),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_output_pipe_3306_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_output_pipe_3306_inst_req_0;
      RPIPE_output_pipe_3306_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_output_pipe_3306_inst_req_1;
      RPIPE_output_pipe_3306_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      output_data_read_3307 <= data_out(15 downto 0);
      output_pipe_read_1_gI: SplitGuardInterface generic map(name => "output_pipe_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      output_pipe_read_1: InputPortRevised -- 
        generic map ( name => "output_pipe_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => output_pipe_pipe_read_req(0),
          oack => output_pipe_pipe_read_ack(0),
          odata => output_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_input_done_pipe_3669_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_3669_inst_req_0;
      WPIPE_input_done_pipe_3669_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_3669_inst_req_1;
      WPIPE_input_done_pipe_3669_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_3670_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendModule_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_1601_start: Boolean;
  signal timer_CP_1601_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_515_inst_req_1 : boolean;
  signal WPIPE_timer_req_515_inst_ack_1 : boolean;
  signal WPIPE_timer_req_515_inst_ack_0 : boolean;
  signal WPIPE_timer_req_515_inst_req_0 : boolean;
  signal RPIPE_timer_resp_520_inst_req_0 : boolean;
  signal RPIPE_timer_resp_520_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_520_inst_req_1 : boolean;
  signal RPIPE_timer_resp_520_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_1601_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1601_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_1601_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1601_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_1601: Block -- control-path 
    signal timer_CP_1601_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_1601_elements(0) <= timer_CP_1601_start;
    timer_CP_1601_symbol <= timer_CP_1601_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/$entry
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_sample_start_
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Sample/req
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Sample/rr
      -- 
    rr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1601_elements(0), ack => RPIPE_timer_resp_520_inst_req_0); -- 
    req_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1601_elements(0), ack => WPIPE_timer_req_515_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Update/$entry
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Update/req
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_update_start_
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Sample/ack
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_sample_completed_
      -- 
    ack_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_515_inst_ack_0, ack => timer_CP_1601_elements(1)); -- 
    req_1619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1601_elements(1), ack => WPIPE_timer_req_515_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Update/$exit
      -- CP-element group 2: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Update/ack
      -- CP-element group 2: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_update_completed_
      -- 
    ack_1620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_515_inst_ack_1, ack => timer_CP_1601_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_update_start_
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_sample_completed_
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Sample/ra
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Update/$entry
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Update/cr
      -- 
    ra_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_520_inst_ack_0, ack => timer_CP_1601_elements(3)); -- 
    cr_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1601_elements(3), ack => RPIPE_timer_resp_520_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_update_completed_
      -- CP-element group 4: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Update/$exit
      -- CP-element group 4: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Update/ca
      -- 
    ca_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_520_inst_ack_1, ack => timer_CP_1601_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_518_to_assign_stmt_521/$exit
      -- CP-element group 5: 	 $exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_1601_elements(2) & timer_CP_1601_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_1601_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_517_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_517_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_520_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_520_inst_req_0;
      RPIPE_timer_resp_520_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_520_inst_req_1;
      RPIPE_timer_resp_520_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_515_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_515_inst_req_0;
      WPIPE_timer_req_515_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_515_inst_req_1;
      WPIPE_timer_req_515_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_517_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_10352_start: Boolean;
  signal timerDaemon_CP_10352_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_resp_3979_inst_req_1 : boolean;
  signal WPIPE_timer_resp_3979_inst_req_0 : boolean;
  signal do_while_stmt_3962_branch_ack_1 : boolean;
  signal phi_stmt_3964_req_0 : boolean;
  signal WPIPE_timer_resp_3979_inst_ack_0 : boolean;
  signal nCOUNTER_3977_3968_buf_req_1 : boolean;
  signal nCOUNTER_3977_3968_buf_req_0 : boolean;
  signal nCOUNTER_3977_3968_buf_ack_1 : boolean;
  signal phi_stmt_3964_req_1 : boolean;
  signal do_while_stmt_3962_branch_ack_0 : boolean;
  signal WPIPE_timer_resp_3979_inst_ack_1 : boolean;
  signal do_while_stmt_3962_branch_req_0 : boolean;
  signal nCOUNTER_3977_3968_buf_ack_0 : boolean;
  signal RPIPE_timer_req_3971_inst_ack_1 : boolean;
  signal RPIPE_timer_req_3971_inst_req_1 : boolean;
  signal RPIPE_timer_req_3971_inst_ack_0 : boolean;
  signal phi_stmt_3964_ack_0 : boolean;
  signal RPIPE_timer_req_3971_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_10352_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_10352_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_10352_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_10352_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_10352: Block -- control-path 
    signal timerDaemon_CP_10352_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_10352_elements(0) <= timerDaemon_CP_10352_start;
    timerDaemon_CP_10352_symbol <= timerDaemon_CP_10352_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_3961/branch_block_stmt_3961__entry__
      -- CP-element group 0: 	 branch_block_stmt_3961/$entry
      -- CP-element group 0: 	 branch_block_stmt_3961/do_while_stmt_3962__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_3961/do_while_stmt_3962__exit__
      -- CP-element group 1: 	 branch_block_stmt_3961/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_3961/branch_block_stmt_3961__exit__
      -- 
    timerDaemon_CP_10352_elements(1) <= timerDaemon_CP_10352_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962__entry__
      -- CP-element group 2: 	 branch_block_stmt_3961/do_while_stmt_3962/$entry
      -- 
    timerDaemon_CP_10352_elements(2) <= timerDaemon_CP_10352_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962__exit__
      -- 
    -- Element group timerDaemon_CP_10352_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_3961/do_while_stmt_3962/loop_back
      -- 
    -- Element group timerDaemon_CP_10352_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_3961/do_while_stmt_3962/condition_done
      -- CP-element group 5: 	 branch_block_stmt_3961/do_while_stmt_3962/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_3961/do_while_stmt_3962/loop_exit/$entry
      -- 
    timerDaemon_CP_10352_elements(5) <= timerDaemon_CP_10352_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_3961/do_while_stmt_3962/loop_body_done
      -- 
    timerDaemon_CP_10352_elements(6) <= timerDaemon_CP_10352_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_10352_elements(7) <= timerDaemon_CP_10352_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_10352_elements(8) <= timerDaemon_CP_10352_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3969_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/loop_body_start
      -- 
    -- Element group timerDaemon_CP_10352_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	40 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/condition_evaluated
      -- 
    condition_evaluated_10376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_10376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10352_elements(10), ack => do_while_stmt_3962_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(14) & timerDaemon_CP_10352_elements(40);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/aggregated_phi_sample_req
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(9) & timerDaemon_CP_10352_elements(15) & timerDaemon_CP_10352_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3969_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/aggregated_phi_sample_ack
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(17) & timerDaemon_CP_10352_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/aggregated_phi_update_req
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(16) & timerDaemon_CP_10352_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(18) & timerDaemon_CP_10352_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(9) & timerDaemon_CP_10352_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(9) & timerDaemon_CP_10352_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_10352_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_update_completed_
      -- 
    -- Element group timerDaemon_CP_10352_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_loopback_trigger
      -- 
    timerDaemon_CP_10352_elements(19) <= timerDaemon_CP_10352_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_loopback_sample_req
      -- 
    phi_stmt_3964_loopback_sample_req_10391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3964_loopback_sample_req_10391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10352_elements(20), ack => phi_stmt_3964_req_1); -- 
    -- Element group timerDaemon_CP_10352_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_entry_trigger
      -- 
    timerDaemon_CP_10352_elements(21) <= timerDaemon_CP_10352_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_entry_sample_req
      -- 
    phi_stmt_3964_entry_sample_req_10394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3964_entry_sample_req_10394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10352_elements(22), ack => phi_stmt_3964_req_0); -- 
    -- Element group timerDaemon_CP_10352_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3964_phi_mux_ack
      -- 
    phi_stmt_3964_phi_mux_ack_10397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3964_ack_0, ack => timerDaemon_CP_10352_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/type_cast_3967_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/type_cast_3967_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/type_cast_3967_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/type_cast_3967_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_10352_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/type_cast_3967_update_start_
      -- CP-element group 25: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/type_cast_3967_update_start__ps
      -- 
    -- Element group timerDaemon_CP_10352_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/type_cast_3967_update_completed__ps
      -- 
    timerDaemon_CP_10352_elements(26) <= timerDaemon_CP_10352_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/type_cast_3967_update_completed_
      -- 
    -- Element group timerDaemon_CP_10352_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_10352_elements(25), ack => timerDaemon_CP_10352_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_sample_start__ps
      -- 
    req_10418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10352_elements(28), ack => nCOUNTER_3977_3968_buf_req_0); -- 
    -- Element group timerDaemon_CP_10352_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_Update/req
      -- CP-element group 29: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_update_start_
      -- CP-element group 29: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_update_start__ps
      -- 
    req_10423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10352_elements(29), ack => nCOUNTER_3977_3968_buf_req_1); -- 
    -- Element group timerDaemon_CP_10352_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_sample_completed__ps
      -- 
    ack_10419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_3977_3968_buf_ack_0, ack => timerDaemon_CP_10352_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/R_nCOUNTER_3968_update_completed__ps
      -- 
    ack_10424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_3977_3968_buf_ack_1, ack => timerDaemon_CP_10352_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3969_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(9) & timerDaemon_CP_10352_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_Sample/rr
      -- 
    rr_10437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10352_elements(33), ack => RPIPE_timer_req_3971_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(11) & timerDaemon_CP_10352_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_update_start_
      -- CP-element group 34: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_Update/$entry
      -- 
    cr_10442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10352_elements(34), ack => RPIPE_timer_req_3971_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(13) & timerDaemon_CP_10352_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_Sample/ra
      -- 
    ra_10438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_3971_inst_ack_0, ack => timerDaemon_CP_10352_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/phi_stmt_3969_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/RPIPE_timer_req_3971_Update/$exit
      -- 
    ca_10443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_3971_inst_ack_1, ack => timerDaemon_CP_10352_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_sample_start_
      -- 
    req_10451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10352_elements(37), ack => WPIPE_timer_resp_3979_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(18) & timerDaemon_CP_10352_elements(36) & timerDaemon_CP_10352_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_Update/req
      -- CP-element group 38: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_update_start_
      -- CP-element group 38: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_Sample/$exit
      -- 
    ack_10452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_3979_inst_ack_0, ack => timerDaemon_CP_10352_elements(38)); -- 
    req_10456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_10352_elements(38), ack => WPIPE_timer_resp_3979_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/WPIPE_timer_resp_3979_Update/ack
      -- 
    ack_10457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_3979_inst_ack_1, ack => timerDaemon_CP_10352_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_10352_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_10352_elements(9), ack => timerDaemon_CP_10352_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_3961/do_while_stmt_3962/do_while_stmt_3962_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_10352_elements(12) & timerDaemon_CP_10352_elements(39);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_10352_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_3961/do_while_stmt_3962/loop_exit/ack
      -- CP-element group 42: 	 branch_block_stmt_3961/do_while_stmt_3962/loop_exit/$exit
      -- 
    ack_10462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3962_branch_ack_0, ack => timerDaemon_CP_10352_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_3961/do_while_stmt_3962/loop_taken/ack
      -- CP-element group 43: 	 branch_block_stmt_3961/do_while_stmt_3962/loop_taken/$exit
      -- 
    ack_10466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3962_branch_ack_1, ack => timerDaemon_CP_10352_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_3961/do_while_stmt_3962/$exit
      -- 
    timerDaemon_CP_10352_elements(44) <= timerDaemon_CP_10352_elements(3);
    timerDaemon_do_while_stmt_3962_terminator_10467: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_3962_terminator_10467", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_10352_elements(6),loop_continue => timerDaemon_CP_10352_elements(43),loop_terminate => timerDaemon_CP_10352_elements(42),loop_back => timerDaemon_CP_10352_elements(4),loop_exit => timerDaemon_CP_10352_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_3964_phi_seq_10425_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_10352_elements(21);
      timerDaemon_CP_10352_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_10352_elements(24);
      timerDaemon_CP_10352_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_10352_elements(26);
      timerDaemon_CP_10352_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_10352_elements(19);
      timerDaemon_CP_10352_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_10352_elements(30);
      timerDaemon_CP_10352_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_10352_elements(31);
      timerDaemon_CP_10352_elements(20) <= phi_mux_reqs(1);
      phi_stmt_3964_phi_seq_10425 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_3964_phi_seq_10425") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_10352_elements(11), 
          phi_sample_ack => timerDaemon_CP_10352_elements(17), 
          phi_update_req => timerDaemon_CP_10352_elements(13), 
          phi_update_ack => timerDaemon_CP_10352_elements(18), 
          phi_mux_ack => timerDaemon_CP_10352_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_10377_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_10352_elements(7);
        preds(1)  <= timerDaemon_CP_10352_elements(8);
        entry_tmerge_10377 : transition_merge -- 
          generic map(name => " entry_tmerge_10377")
          port map (preds => preds, symbol_out => timerDaemon_CP_10352_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_3964 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_3971_wire : std_logic_vector(0 downto 0);
    signal konst_3975_wire_constant : std_logic_vector(63 downto 0);
    signal konst_3983_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_3977 : std_logic_vector(63 downto 0);
    signal nCOUNTER_3977_3968_buffered : std_logic_vector(63 downto 0);
    signal req_3969 : std_logic_vector(0 downto 0);
    signal type_cast_3967_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_3975_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_3983_wire_constant <= "1";
    type_cast_3967_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_3964: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3967_wire_constant & nCOUNTER_3977_3968_buffered;
      req <= phi_stmt_3964_req_0 & phi_stmt_3964_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3964",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3964_ack_0,
          idata => idata,
          odata => COUNTER_3964,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3964
    nCOUNTER_3977_3968_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_3977_3968_buf_req_0;
      nCOUNTER_3977_3968_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_3977_3968_buf_req_1;
      nCOUNTER_3977_3968_buf_ack_1<= rack(0);
      nCOUNTER_3977_3968_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_3977_3968_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_3977,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_3977_3968_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_3969
    process(RPIPE_timer_req_3971_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_3971_wire(0 downto 0);
      req_3969 <= tmp_var; -- 
    end process;
    do_while_stmt_3962_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_3983_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_3962_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_3962_branch_req_0,
          ack0 => do_while_stmt_3962_branch_ack_0,
          ack1 => do_while_stmt_3962_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_3976_inst
    process(COUNTER_3964) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_3964, konst_3975_wire_constant, tmp_var);
      nCOUNTER_3977 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_3971_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_3971_inst_req_0;
      RPIPE_timer_req_3971_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_3971_inst_req_1;
      RPIPE_timer_req_3971_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_3971_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_3979_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_3979_inst_req_0;
      WPIPE_timer_resp_3979_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_3979_inst_req_1;
      WPIPE_timer_resp_3979_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_3969(0);
      data_in <= COUNTER_3964;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(27 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(37 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(127 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(7 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(7 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(7 downto 0);
      input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_row_in :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(47 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(47 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(47 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(79 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      sendB_call_reqs : out  std_logic_vector(0 downto 0);
      sendB_call_acks : in   std_logic_vector(0 downto 0);
      sendB_call_data : out  std_logic_vector(31 downto 0);
      sendB_call_tag  :  out  std_logic_vector(0 downto 0);
      sendB_return_reqs : out  std_logic_vector(0 downto 0);
      sendB_return_acks : in   std_logic_vector(0 downto 0);
      sendB_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_data : in   std_logic_vector(7 downto 0);
      input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_data : in   std_logic_vector(7 downto 0);
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_data : in   std_logic_vector(7 downto 0);
      input_pipe4_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(7 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(7 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(7 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_num_chl :  std_logic_vector(15 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(79 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(79 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendB
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendB
  signal sendB_size :  std_logic_vector(31 downto 0);
  signal sendB_in_args    : std_logic_vector(31 downto 0);
  signal sendB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendB_tag_out   : std_logic_vector(1 downto 0);
  signal sendB_start_req : std_logic;
  signal sendB_start_ack : std_logic;
  signal sendB_fin_req   : std_logic;
  signal sendB_fin_ack : std_logic;
  -- caller side aggregated signals for module sendB
  signal sendB_call_reqs: std_logic_vector(0 downto 0);
  signal sendB_call_acks: std_logic_vector(0 downto 0);
  signal sendB_return_reqs: std_logic_vector(0 downto 0);
  signal sendB_return_acks: std_logic_vector(0 downto 0);
  signal sendB_call_data: std_logic_vector(31 downto 0);
  signal sendB_call_tag: std_logic_vector(0 downto 0);
  signal sendB_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendModule
  component sendModule is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      output_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
      output_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
      output_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendModule
  signal sendModule_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendModule_tag_out   : std_logic_vector(1 downto 0);
  signal sendModule_start_req : std_logic;
  signal sendModule_start_ack : std_logic;
  signal sendModule_fin_req   : std_logic;
  signal sendModule_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(7 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(7 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe2
  signal input_pipe2_pipe_write_data: std_logic_vector(7 downto 0);
  signal input_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe2
  signal input_pipe2_pipe_read_data: std_logic_vector(7 downto 0);
  signal input_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe3
  signal input_pipe3_pipe_write_data: std_logic_vector(7 downto 0);
  signal input_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe3
  signal input_pipe3_pipe_read_data: std_logic_vector(7 downto 0);
  signal input_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe4
  signal input_pipe4_pipe_write_data: std_logic_vector(7 downto 0);
  signal input_pipe4_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe4
  signal input_pipe4_pipe_read_data: std_logic_vector(7 downto 0);
  signal input_pipe4_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(7 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(7 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe2
  signal kernel_pipe2_pipe_write_data: std_logic_vector(7 downto 0);
  signal kernel_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe2
  signal kernel_pipe2_pipe_read_data: std_logic_vector(7 downto 0);
  signal kernel_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe3
  signal kernel_pipe3_pipe_write_data: std_logic_vector(7 downto 0);
  signal kernel_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe3
  signal kernel_pipe3_pipe_read_data: std_logic_vector(7 downto 0);
  signal kernel_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe output_pipe
  signal output_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe output_pipe
  signal output_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal output_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal output_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_row_in <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 48,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      row_in => access_T_row_in,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(20 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 0),
      input_pipe2_pipe_write_req => input_pipe2_pipe_write_req(0 downto 0),
      input_pipe2_pipe_write_ack => input_pipe2_pipe_write_ack(0 downto 0),
      input_pipe2_pipe_write_data => input_pipe2_pipe_write_data(7 downto 0),
      input_pipe3_pipe_write_req => input_pipe3_pipe_write_req(0 downto 0),
      input_pipe3_pipe_write_ack => input_pipe3_pipe_write_ack(0 downto 0),
      input_pipe3_pipe_write_data => input_pipe3_pipe_write_data(7 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(7 downto 0),
      input_pipe4_pipe_write_req => input_pipe4_pipe_write_req(0 downto 0),
      input_pipe4_pipe_write_ack => input_pipe4_pipe_write_ack(0 downto 0),
      input_pipe4_pipe_write_data => input_pipe4_pipe_write_data(7 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(20 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(7 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      output_pipe_pipe_write_req => output_pipe_pipe_write_req(1 downto 1),
      output_pipe_pipe_write_ack => output_pipe_pipe_write_ack(1 downto 1),
      output_pipe_pipe_write_data => output_pipe_pipe_write_data(31 downto 16),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(47 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(79 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      sendB_call_reqs => sendB_call_reqs(0 downto 0),
      sendB_call_acks => sendB_call_acks(0 downto 0),
      sendB_call_data => sendB_call_data(31 downto 0),
      sendB_call_tag => sendB_call_tag(0 downto 0),
      sendB_return_reqs => sendB_return_reqs(0 downto 0),
      sendB_return_acks => sendB_return_acks(0 downto 0),
      sendB_return_tag => sendB_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe2_pipe_read_req => input_pipe2_pipe_read_req(0 downto 0),
      input_pipe2_pipe_read_ack => input_pipe2_pipe_read_ack(0 downto 0),
      input_pipe2_pipe_read_data => input_pipe2_pipe_read_data(7 downto 0),
      input_pipe3_pipe_read_req => input_pipe3_pipe_read_req(0 downto 0),
      input_pipe3_pipe_read_ack => input_pipe3_pipe_read_ack(0 downto 0),
      input_pipe3_pipe_read_data => input_pipe3_pipe_read_data(7 downto 0),
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(7 downto 0),
      kernel_pipe2_pipe_read_req => kernel_pipe2_pipe_read_req(0 downto 0),
      kernel_pipe2_pipe_read_ack => kernel_pipe2_pipe_read_ack(0 downto 0),
      kernel_pipe2_pipe_read_data => kernel_pipe2_pipe_read_data(7 downto 0),
      kernel_pipe3_pipe_read_req => kernel_pipe3_pipe_read_req(0 downto 0),
      kernel_pipe3_pipe_read_ack => kernel_pipe3_pipe_read_ack(0 downto 0),
      kernel_pipe3_pipe_read_data => kernel_pipe3_pipe_read_data(7 downto 0),
      input_pipe4_pipe_read_req => input_pipe4_pipe_read_req(0 downto 0),
      input_pipe4_pipe_read_ack => input_pipe4_pipe_read_ack(0 downto 0),
      input_pipe4_pipe_read_data => input_pipe4_pipe_read_data(7 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(7 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(1 downto 1),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(1 downto 1),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(15 downto 8),
      output_pipe_pipe_write_req => output_pipe_pipe_write_req(0 downto 0),
      output_pipe_pipe_write_ack => output_pipe_pipe_write_ack(0 downto 0),
      output_pipe_pipe_write_data => output_pipe_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(79 downto 16);
  loadKernelChannel_num_chl <= loadKernelChannel_in_args(15 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 80,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      num_chl => loadKernelChannel_num_chl,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(1 downto 1),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(1 downto 1),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(15 downto 8),
      kernel_pipe2_pipe_write_req => kernel_pipe2_pipe_write_req(0 downto 0),
      kernel_pipe2_pipe_write_ack => kernel_pipe2_pipe_write_ack(0 downto 0),
      kernel_pipe2_pipe_write_data => kernel_pipe2_pipe_write_data(7 downto 0),
      kernel_pipe3_pipe_write_req => kernel_pipe3_pipe_write_req(0 downto 0),
      kernel_pipe3_pipe_write_ack => kernel_pipe3_pipe_write_ack(0 downto 0),
      kernel_pipe3_pipe_write_data => kernel_pipe3_pipe_write_data(7 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(7 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(15 downto 0),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module sendB
  sendB_size <= sendB_in_args(31 downto 0);
  -- call arbiter for module sendB
  sendB_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendB_call_reqs,
      call_acks => sendB_call_acks,
      return_reqs => sendB_return_reqs,
      return_acks => sendB_return_acks,
      call_data  => sendB_call_data,
      call_tag  => sendB_call_tag,
      return_tag  => sendB_return_tag,
      call_mtag => sendB_tag_in,
      return_mtag => sendB_tag_out,
      call_mreq => sendB_start_req,
      call_mack => sendB_start_ack,
      return_mreq => sendB_fin_req,
      return_mack => sendB_fin_ack,
      call_mdata => sendB_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendB_instance:sendB-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendB_size,
      start_req => sendB_start_req,
      start_ack => sendB_start_ack,
      fin_req => sendB_fin_req,
      fin_ack => sendB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(37 downto 19),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 2),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      tag_in => sendB_tag_in,
      tag_out => sendB_tag_out-- 
    ); -- 
  -- module sendModule
  sendModule_instance:sendModule-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendModule_start_req,
      start_ack => sendModule_start_ack,
      fin_req => sendModule_fin_req,
      fin_ack => sendModule_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      output_pipe_pipe_read_req => output_pipe_pipe_read_req(1 downto 0),
      output_pipe_pipe_read_ack => output_pipe_pipe_read_ack(1 downto 0),
      output_pipe_pipe_read_data => output_pipe_pipe_read_data(31 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(7 downto 0),
      tag_in => sendModule_tag_in,
      tag_out => sendModule_tag_out-- 
    ); -- 
  -- module will be run forever 
  sendModule_tag_in <= (others => '0');
  sendModule_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => sendModule_start_req, start_ack => sendModule_start_ack,  fin_req => sendModule_fin_req,  fin_ack => sendModule_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 2,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe2_pipe_read_req,
      read_ack => input_pipe2_pipe_read_ack,
      read_data => input_pipe2_pipe_read_data,
      write_req => input_pipe2_pipe_write_req,
      write_ack => input_pipe2_pipe_write_ack,
      write_data => input_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe3_pipe_read_req,
      read_ack => input_pipe3_pipe_read_ack,
      read_data => input_pipe3_pipe_read_data,
      write_req => input_pipe3_pipe_write_req,
      write_ack => input_pipe3_pipe_write_ack,
      write_data => input_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe4",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe4_pipe_read_req,
      read_ack => input_pipe4_pipe_read_ack,
      read_data => input_pipe4_pipe_read_data,
      write_req => input_pipe4_pipe_write_req,
      write_ack => input_pipe4_pipe_write_ack,
      write_data => input_pipe4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe2_pipe_read_req,
      read_ack => kernel_pipe2_pipe_read_ack,
      read_data => kernel_pipe2_pipe_read_data,
      write_req => kernel_pipe2_pipe_write_req,
      write_ack => kernel_pipe2_pipe_write_ack,
      write_data => kernel_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe3_pipe_read_req,
      read_ack => kernel_pipe3_pipe_read_ack,
      read_data => kernel_pipe3_pipe_read_data,
      write_req => kernel_pipe3_pipe_write_req,
      write_ack => kernel_pipe3_pipe_write_ack,
      write_data => kernel_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe output_pipe",
      num_reads => 2,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 10 --
    )
    port map( -- 
      read_req => output_pipe_pipe_read_req,
      read_ack => output_pipe_pipe_read_ack,
      read_data => output_pipe_pipe_read_data,
      write_req => output_pipe_pipe_write_req,
      write_ack => output_pipe_pipe_write_ack,
      write_data => output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 11 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
