-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ct_core is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(9 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity ct_core;
architecture ct_core_arch of ct_core is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ct_core_CP_34_start: Boolean;
  signal ct_core_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_ConvTranspose_input_pipe_517_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_706_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_688_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_ack_0 : boolean;
  signal type_cast_485_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_688_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_req_1 : boolean;
  signal type_cast_45_inst_req_0 : boolean;
  signal type_cast_45_inst_ack_0 : boolean;
  signal type_cast_45_inst_req_1 : boolean;
  signal type_cast_539_inst_ack_0 : boolean;
  signal type_cast_45_inst_ack_1 : boolean;
  signal array_obj_ref_464_index_offset_ack_1 : boolean;
  signal array_obj_ref_464_index_offset_req_1 : boolean;
  signal type_cast_485_inst_ack_1 : boolean;
  signal array_obj_ref_464_index_offset_ack_0 : boolean;
  signal array_obj_ref_464_index_offset_req_0 : boolean;
  signal type_cast_485_inst_req_1 : boolean;
  signal type_cast_485_inst_ack_0 : boolean;
  signal type_cast_539_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_27_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_27_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_27_inst_req_1 : boolean;
  signal type_cast_539_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_27_inst_ack_1 : boolean;
  signal type_cast_1388_inst_req_0 : boolean;
  signal ptr_deref_601_store_0_ack_1 : boolean;
  signal type_cast_32_inst_req_0 : boolean;
  signal type_cast_32_inst_ack_0 : boolean;
  signal type_cast_32_inst_req_1 : boolean;
  signal type_cast_32_inst_ack_1 : boolean;
  signal ptr_deref_1018_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_41_inst_ack_1 : boolean;
  signal array_obj_ref_671_index_offset_ack_1 : boolean;
  signal array_obj_ref_671_index_offset_req_1 : boolean;
  signal addr_of_672_final_reg_ack_1 : boolean;
  signal type_cast_692_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_ack_0 : boolean;
  signal type_cast_472_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_141_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_481_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_0 : boolean;
  signal add_dest_dim0_init_946_972_buf_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_481_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_1 : boolean;
  signal type_cast_539_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 : boolean;
  signal array_obj_ref_671_index_offset_ack_0 : boolean;
  signal ptr_deref_601_store_0_req_1 : boolean;
  signal addr_of_672_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_481_inst_req_0 : boolean;
  signal type_cast_57_inst_req_0 : boolean;
  signal next_add_src_1111_981_buf_req_1 : boolean;
  signal type_cast_57_inst_ack_0 : boolean;
  signal type_cast_57_inst_req_1 : boolean;
  signal type_cast_57_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_66_inst_ack_1 : boolean;
  signal W_ov_1028_delayed_6_0_1028_inst_req_1 : boolean;
  signal type_cast_1368_inst_req_1 : boolean;
  signal array_obj_ref_671_index_offset_req_0 : boolean;
  signal add_dest_dim0_init_946_972_buf_req_0 : boolean;
  signal type_cast_1418_inst_ack_1 : boolean;
  signal type_cast_70_inst_req_0 : boolean;
  signal type_cast_70_inst_ack_0 : boolean;
  signal type_cast_70_inst_req_1 : boolean;
  signal type_cast_70_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_675_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_481_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_ack_1 : boolean;
  signal type_cast_1378_inst_ack_1 : boolean;
  signal type_cast_82_inst_req_0 : boolean;
  signal type_cast_82_inst_ack_0 : boolean;
  signal type_cast_82_inst_req_1 : boolean;
  signal type_cast_82_inst_ack_1 : boolean;
  signal phi_stmt_974_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_91_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_req_0 : boolean;
  signal type_cast_95_inst_req_0 : boolean;
  signal type_cast_95_inst_ack_0 : boolean;
  signal type_cast_95_inst_req_1 : boolean;
  signal type_cast_95_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_675_inst_req_1 : boolean;
  signal next_add_src_1111_981_buf_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_req_1 : boolean;
  signal next_add_src_1111_981_buf_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_ack_1 : boolean;
  signal type_cast_679_inst_ack_1 : boolean;
  signal type_cast_503_inst_ack_1 : boolean;
  signal type_cast_107_inst_req_0 : boolean;
  signal type_cast_107_inst_ack_0 : boolean;
  signal type_cast_107_inst_req_1 : boolean;
  signal type_cast_107_inst_ack_1 : boolean;
  signal next_input_dim1_1143_965_buf_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_req_1 : boolean;
  signal add_dest_dim0_init_946_972_buf_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_116_inst_ack_1 : boolean;
  signal type_cast_679_inst_req_1 : boolean;
  signal next_input_dim2_1133_969_buf_req_1 : boolean;
  signal ptr_deref_601_store_0_ack_0 : boolean;
  signal addr_of_672_final_reg_ack_0 : boolean;
  signal type_cast_503_inst_req_1 : boolean;
  signal type_cast_120_inst_req_0 : boolean;
  signal type_cast_120_inst_ack_0 : boolean;
  signal type_cast_120_inst_req_1 : boolean;
  signal type_cast_120_inst_ack_1 : boolean;
  signal type_cast_692_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 : boolean;
  signal if_stmt_615_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_1 : boolean;
  signal next_input_dim1_1143_965_buf_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 : boolean;
  signal ptr_deref_601_store_0_req_0 : boolean;
  signal type_cast_132_inst_req_0 : boolean;
  signal type_cast_132_inst_ack_0 : boolean;
  signal type_cast_132_inst_req_1 : boolean;
  signal type_cast_132_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 : boolean;
  signal addr_of_465_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 : boolean;
  signal type_cast_642_inst_ack_0 : boolean;
  signal type_cast_642_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_589_inst_ack_1 : boolean;
  signal type_cast_593_inst_ack_1 : boolean;
  signal type_cast_320_inst_req_0 : boolean;
  signal type_cast_320_inst_ack_0 : boolean;
  signal type_cast_320_inst_req_1 : boolean;
  signal type_cast_320_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_688_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_req_0 : boolean;
  signal type_cast_593_inst_req_1 : boolean;
  signal addr_of_672_final_reg_req_0 : boolean;
  signal type_cast_557_inst_ack_1 : boolean;
  signal type_cast_503_inst_ack_0 : boolean;
  signal type_cast_145_inst_req_0 : boolean;
  signal type_cast_145_inst_ack_0 : boolean;
  signal type_cast_145_inst_req_1 : boolean;
  signal type_cast_145_inst_ack_1 : boolean;
  signal W_ov_1028_delayed_6_0_1028_inst_ack_1 : boolean;
  signal type_cast_472_inst_req_1 : boolean;
  signal type_cast_557_inst_req_1 : boolean;
  signal type_cast_575_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_ack_1 : boolean;
  signal type_cast_157_inst_req_0 : boolean;
  signal type_cast_157_inst_ack_0 : boolean;
  signal type_cast_157_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_ack_0 : boolean;
  signal type_cast_157_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_675_inst_ack_0 : boolean;
  signal type_cast_575_inst_req_1 : boolean;
  signal if_stmt_615_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_ack_0 : boolean;
  signal type_cast_472_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_535_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_166_inst_ack_1 : boolean;
  signal type_cast_557_inst_ack_0 : boolean;
  signal type_cast_170_inst_req_0 : boolean;
  signal type_cast_1378_inst_ack_0 : boolean;
  signal type_cast_170_inst_ack_0 : boolean;
  signal type_cast_170_inst_req_1 : boolean;
  signal type_cast_170_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_675_inst_req_0 : boolean;
  signal type_cast_692_inst_ack_0 : boolean;
  signal type_cast_472_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_ack_1 : boolean;
  signal type_cast_679_inst_ack_0 : boolean;
  signal type_cast_557_inst_req_0 : boolean;
  signal type_cast_503_inst_req_0 : boolean;
  signal type_cast_182_inst_req_0 : boolean;
  signal type_cast_182_inst_ack_0 : boolean;
  signal type_cast_182_inst_req_1 : boolean;
  signal type_cast_182_inst_ack_1 : boolean;
  signal type_cast_692_inst_req_0 : boolean;
  signal next_add_src_1111_981_buf_ack_0 : boolean;
  signal type_cast_575_inst_ack_0 : boolean;
  signal type_cast_575_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_191_inst_ack_1 : boolean;
  signal type_cast_679_inst_req_0 : boolean;
  signal type_cast_195_inst_req_0 : boolean;
  signal type_cast_195_inst_ack_0 : boolean;
  signal type_cast_195_inst_req_1 : boolean;
  signal type_cast_195_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_ack_1 : boolean;
  signal add_dest_dim0_init_946_972_buf_ack_0 : boolean;
  signal type_cast_207_inst_req_0 : boolean;
  signal type_cast_207_inst_ack_0 : boolean;
  signal type_cast_207_inst_req_1 : boolean;
  signal next_input_dim1_1143_965_buf_ack_1 : boolean;
  signal type_cast_207_inst_ack_1 : boolean;
  signal if_stmt_615_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_216_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_216_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_216_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_216_inst_ack_1 : boolean;
  signal phi_stmt_881_req_0 : boolean;
  signal type_cast_220_inst_req_0 : boolean;
  signal type_cast_220_inst_ack_0 : boolean;
  signal type_cast_220_inst_req_1 : boolean;
  signal type_cast_220_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_228_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_228_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_468_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_228_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_228_inst_ack_1 : boolean;
  signal type_cast_232_inst_req_0 : boolean;
  signal type_cast_232_inst_ack_0 : boolean;
  signal type_cast_232_inst_req_1 : boolean;
  signal type_cast_232_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_468_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_241_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_241_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_241_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_241_inst_ack_1 : boolean;
  signal type_cast_245_inst_req_0 : boolean;
  signal type_cast_521_inst_ack_1 : boolean;
  signal type_cast_245_inst_ack_0 : boolean;
  signal type_cast_245_inst_req_1 : boolean;
  signal type_cast_245_inst_ack_1 : boolean;
  signal type_cast_665_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_253_inst_req_0 : boolean;
  signal type_cast_521_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_253_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_468_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_253_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_253_inst_ack_1 : boolean;
  signal ptr_deref_1018_load_0_req_0 : boolean;
  signal type_cast_257_inst_req_0 : boolean;
  signal type_cast_257_inst_ack_0 : boolean;
  signal type_cast_257_inst_req_1 : boolean;
  signal type_cast_257_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_468_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_266_inst_req_0 : boolean;
  signal type_cast_521_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_266_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_266_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_266_inst_ack_1 : boolean;
  signal type_cast_1428_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_req_1 : boolean;
  signal type_cast_270_inst_req_0 : boolean;
  signal type_cast_521_inst_req_0 : boolean;
  signal type_cast_270_inst_ack_0 : boolean;
  signal type_cast_270_inst_req_1 : boolean;
  signal type_cast_1378_inst_req_0 : boolean;
  signal type_cast_270_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_278_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_278_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_278_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_278_inst_ack_1 : boolean;
  signal phi_stmt_881_req_1 : boolean;
  signal type_cast_282_inst_req_0 : boolean;
  signal type_cast_282_inst_ack_0 : boolean;
  signal type_cast_282_inst_req_1 : boolean;
  signal type_cast_282_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_ack_1 : boolean;
  signal type_cast_1418_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_ack_1 : boolean;
  signal type_cast_642_inst_ack_1 : boolean;
  signal type_cast_642_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_553_inst_req_1 : boolean;
  signal type_cast_295_inst_req_0 : boolean;
  signal type_cast_295_inst_ack_0 : boolean;
  signal type_cast_295_inst_req_1 : boolean;
  signal type_cast_295_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_303_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_303_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_303_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_303_inst_ack_1 : boolean;
  signal type_cast_307_inst_req_0 : boolean;
  signal type_cast_307_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_571_inst_req_1 : boolean;
  signal type_cast_307_inst_req_1 : boolean;
  signal type_cast_307_inst_ack_1 : boolean;
  signal addr_of_465_final_reg_ack_1 : boolean;
  signal type_cast_330_inst_req_0 : boolean;
  signal type_cast_330_inst_ack_0 : boolean;
  signal type_cast_330_inst_req_1 : boolean;
  signal type_cast_330_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_688_inst_req_1 : boolean;
  signal phi_stmt_978_req_1 : boolean;
  signal type_cast_593_inst_ack_0 : boolean;
  signal type_cast_339_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_ack_0 : boolean;
  signal type_cast_339_inst_ack_0 : boolean;
  signal type_cast_339_inst_req_1 : boolean;
  signal type_cast_339_inst_ack_1 : boolean;
  signal type_cast_593_inst_req_0 : boolean;
  signal type_cast_358_inst_req_0 : boolean;
  signal type_cast_358_inst_ack_0 : boolean;
  signal type_cast_358_inst_req_1 : boolean;
  signal type_cast_358_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_ack_1 : boolean;
  signal type_cast_362_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_req_1 : boolean;
  signal type_cast_362_inst_ack_0 : boolean;
  signal type_cast_362_inst_req_1 : boolean;
  signal type_cast_362_inst_ack_1 : boolean;
  signal next_input_dim2_1133_969_buf_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_req_1 : boolean;
  signal type_cast_371_inst_req_0 : boolean;
  signal type_cast_371_inst_ack_0 : boolean;
  signal addr_of_465_final_reg_ack_0 : boolean;
  signal next_input_dim1_1143_965_buf_req_0 : boolean;
  signal type_cast_371_inst_req_1 : boolean;
  signal type_cast_371_inst_ack_1 : boolean;
  signal addr_of_465_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_499_inst_req_0 : boolean;
  signal type_cast_380_inst_req_0 : boolean;
  signal type_cast_380_inst_ack_0 : boolean;
  signal type_cast_380_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_517_inst_ack_0 : boolean;
  signal type_cast_380_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_req_0 : boolean;
  signal type_cast_1388_inst_ack_1 : boolean;
  signal next_input_dim2_1133_969_buf_req_0 : boolean;
  signal if_stmt_393_branch_req_0 : boolean;
  signal next_input_dim2_1133_969_buf_ack_0 : boolean;
  signal if_stmt_393_branch_ack_1 : boolean;
  signal if_stmt_393_branch_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_req_1 : boolean;
  signal phi_stmt_974_req_1 : boolean;
  signal if_stmt_408_branch_req_0 : boolean;
  signal if_stmt_408_branch_ack_1 : boolean;
  signal if_stmt_408_branch_ack_0 : boolean;
  signal type_cast_435_inst_req_0 : boolean;
  signal type_cast_435_inst_ack_0 : boolean;
  signal type_cast_435_inst_req_1 : boolean;
  signal type_cast_435_inst_ack_1 : boolean;
  signal addr_of_1026_final_reg_ack_1 : boolean;
  signal type_cast_710_inst_req_0 : boolean;
  signal type_cast_710_inst_ack_0 : boolean;
  signal type_cast_710_inst_req_1 : boolean;
  signal type_cast_710_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_724_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0 : boolean;
  signal addr_of_1026_final_reg_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_ack_1 : boolean;
  signal type_cast_728_inst_req_0 : boolean;
  signal type_cast_728_inst_ack_0 : boolean;
  signal type_cast_728_inst_req_1 : boolean;
  signal type_cast_728_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1430_inst_req_0 : boolean;
  signal phi_stmt_970_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_742_inst_ack_1 : boolean;
  signal type_cast_1368_inst_ack_1 : boolean;
  signal type_cast_746_inst_req_0 : boolean;
  signal type_cast_746_inst_ack_0 : boolean;
  signal type_cast_746_inst_req_1 : boolean;
  signal type_cast_746_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_ack_0 : boolean;
  signal phi_stmt_970_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_760_inst_ack_1 : boolean;
  signal W_ov_1028_delayed_6_0_1028_inst_ack_0 : boolean;
  signal type_cast_764_inst_req_0 : boolean;
  signal type_cast_764_inst_ack_0 : boolean;
  signal type_cast_764_inst_req_1 : boolean;
  signal type_cast_764_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_778_inst_ack_1 : boolean;
  signal array_obj_ref_1025_index_offset_ack_1 : boolean;
  signal array_obj_ref_1025_index_offset_req_1 : boolean;
  signal type_cast_782_inst_req_0 : boolean;
  signal type_cast_782_inst_ack_0 : boolean;
  signal type_cast_782_inst_req_1 : boolean;
  signal type_cast_1388_inst_req_1 : boolean;
  signal type_cast_782_inst_ack_1 : boolean;
  signal array_obj_ref_1013_index_offset_ack_1 : boolean;
  signal array_obj_ref_1013_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_ack_0 : boolean;
  signal phi_stmt_970_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_796_inst_ack_1 : boolean;
  signal W_ov_1028_delayed_6_0_1028_inst_req_0 : boolean;
  signal type_cast_800_inst_req_0 : boolean;
  signal type_cast_800_inst_ack_0 : boolean;
  signal type_cast_800_inst_req_1 : boolean;
  signal type_cast_800_inst_ack_1 : boolean;
  signal type_cast_665_inst_ack_0 : boolean;
  signal next_add_dest_dim1_1121_977_buf_ack_1 : boolean;
  signal next_add_dest_dim1_1121_977_buf_req_1 : boolean;
  signal addr_of_1026_final_reg_ack_0 : boolean;
  signal next_add_dest_dim0_1127_973_buf_ack_1 : boolean;
  signal next_add_dest_dim0_1127_973_buf_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_req_0 : boolean;
  signal ptr_deref_808_store_0_req_0 : boolean;
  signal ptr_deref_808_store_0_ack_0 : boolean;
  signal ptr_deref_808_store_0_req_1 : boolean;
  signal next_add_dest_dim1_1121_977_buf_ack_0 : boolean;
  signal ptr_deref_808_store_0_ack_1 : boolean;
  signal array_obj_ref_1025_index_offset_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_ack_0 : boolean;
  signal next_add_dest_dim1_1121_977_buf_req_0 : boolean;
  signal type_cast_1388_inst_ack_0 : boolean;
  signal if_stmt_822_branch_req_0 : boolean;
  signal phi_stmt_978_ack_0 : boolean;
  signal if_stmt_822_branch_ack_1 : boolean;
  signal if_stmt_822_branch_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1430_inst_ack_1 : boolean;
  signal if_stmt_837_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1430_inst_ack_0 : boolean;
  signal phi_stmt_966_ack_0 : boolean;
  signal if_stmt_837_branch_ack_1 : boolean;
  signal if_stmt_837_branch_ack_0 : boolean;
  signal next_add_dest_dim0_1127_973_buf_ack_0 : boolean;
  signal if_stmt_1465_branch_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_req_1 : boolean;
  signal type_cast_864_inst_req_0 : boolean;
  signal type_cast_864_inst_ack_0 : boolean;
  signal type_cast_864_inst_req_1 : boolean;
  signal type_cast_864_inst_ack_1 : boolean;
  signal addr_of_1014_final_reg_ack_1 : boolean;
  signal phi_stmt_966_req_0 : boolean;
  signal addr_of_1026_final_reg_req_0 : boolean;
  signal array_obj_ref_1013_index_offset_ack_0 : boolean;
  signal array_obj_ref_893_index_offset_req_0 : boolean;
  signal array_obj_ref_893_index_offset_ack_0 : boolean;
  signal array_obj_ref_893_index_offset_req_1 : boolean;
  signal array_obj_ref_893_index_offset_ack_1 : boolean;
  signal addr_of_1014_final_reg_req_1 : boolean;
  signal array_obj_ref_1025_index_offset_req_0 : boolean;
  signal phi_stmt_881_ack_0 : boolean;
  signal type_cast_458_inst_req_0 : boolean;
  signal type_cast_1418_inst_req_0 : boolean;
  signal addr_of_894_final_reg_req_0 : boolean;
  signal type_cast_1378_inst_req_1 : boolean;
  signal addr_of_894_final_reg_ack_0 : boolean;
  signal addr_of_894_final_reg_req_1 : boolean;
  signal addr_of_894_final_reg_ack_1 : boolean;
  signal ptr_deref_1018_load_0_ack_1 : boolean;
  signal phi_stmt_452_req_0 : boolean;
  signal ptr_deref_1018_load_0_req_1 : boolean;
  signal type_cast_665_inst_req_1 : boolean;
  signal add_dest_dim1_init_951_976_buf_ack_1 : boolean;
  signal next_add_dest_dim0_1127_973_buf_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1430_inst_req_1 : boolean;
  signal ptr_deref_897_store_0_req_0 : boolean;
  signal add_dest_dim1_init_951_976_buf_req_1 : boolean;
  signal ptr_deref_897_store_0_ack_0 : boolean;
  signal ptr_deref_897_store_0_req_1 : boolean;
  signal ptr_deref_897_store_0_ack_1 : boolean;
  signal add_dest_dim1_init_951_976_buf_ack_0 : boolean;
  signal phi_stmt_978_req_0 : boolean;
  signal if_stmt_912_branch_req_0 : boolean;
  signal add_dest_dim1_init_951_976_buf_req_0 : boolean;
  signal phi_stmt_966_req_1 : boolean;
  signal if_stmt_912_branch_ack_1 : boolean;
  signal if_stmt_912_branch_ack_0 : boolean;
  signal array_obj_ref_1013_index_offset_req_0 : boolean;
  signal if_stmt_1465_branch_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1 : boolean;
  signal type_cast_665_inst_ack_1 : boolean;
  signal call_stmt_923_call_req_0 : boolean;
  signal call_stmt_923_call_ack_0 : boolean;
  signal call_stmt_923_call_req_1 : boolean;
  signal call_stmt_923_call_ack_1 : boolean;
  signal phi_stmt_659_req_1 : boolean;
  signal do_while_stmt_956_branch_req_0 : boolean;
  signal type_cast_1428_inst_req_0 : boolean;
  signal addr_of_1014_final_reg_ack_0 : boolean;
  signal type_cast_1418_inst_ack_0 : boolean;
  signal phi_stmt_958_req_1 : boolean;
  signal phi_stmt_958_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_ack_1 : boolean;
  signal phi_stmt_974_ack_0 : boolean;
  signal phi_stmt_958_ack_0 : boolean;
  signal addr_of_1014_final_reg_req_0 : boolean;
  signal phi_stmt_659_ack_0 : boolean;
  signal type_cast_1428_inst_req_1 : boolean;
  signal type_cast_1428_inst_ack_1 : boolean;
  signal next_input_dim0_1149_961_buf_req_0 : boolean;
  signal next_input_dim0_1149_961_buf_ack_0 : boolean;
  signal next_input_dim0_1149_961_buf_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_req_0 : boolean;
  signal next_input_dim0_1149_961_buf_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0 : boolean;
  signal phi_stmt_962_req_1 : boolean;
  signal phi_stmt_962_req_0 : boolean;
  signal phi_stmt_962_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1439_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1439_inst_req_1 : boolean;
  signal ptr_deref_1032_store_0_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1439_inst_ack_0 : boolean;
  signal ptr_deref_1032_store_0_ack_0 : boolean;
  signal ptr_deref_1032_store_0_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1439_inst_req_0 : boolean;
  signal ptr_deref_1032_store_0_ack_1 : boolean;
  signal phi_stmt_659_req_0 : boolean;
  signal W_dim2_limit_1039_delayed_1_0_1040_inst_req_0 : boolean;
  signal W_dim2_limit_1039_delayed_1_0_1040_inst_ack_0 : boolean;
  signal W_dim2_limit_1039_delayed_1_0_1040_inst_req_1 : boolean;
  signal W_dim2_limit_1039_delayed_1_0_1040_inst_ack_1 : boolean;
  signal SUB_u16_u16_1051_inst_req_0 : boolean;
  signal SUB_u16_u16_1051_inst_ack_0 : boolean;
  signal type_cast_887_inst_ack_1 : boolean;
  signal SUB_u16_u16_1051_inst_req_1 : boolean;
  signal SUB_u16_u16_1051_inst_ack_1 : boolean;
  signal W_nid1_true3_1092_delayed_1_0_1099_inst_req_0 : boolean;
  signal W_nid1_true3_1092_delayed_1_0_1099_inst_ack_0 : boolean;
  signal type_cast_887_inst_req_1 : boolean;
  signal W_nid1_true3_1092_delayed_1_0_1099_inst_req_1 : boolean;
  signal W_nid1_true3_1092_delayed_1_0_1099_inst_ack_1 : boolean;
  signal type_cast_1408_inst_ack_1 : boolean;
  signal type_cast_1368_inst_ack_0 : boolean;
  signal type_cast_1368_inst_req_0 : boolean;
  signal type_cast_1408_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1436_inst_ack_1 : boolean;
  signal type_cast_1408_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1436_inst_req_1 : boolean;
  signal SUB_u16_u16_1153_inst_req_0 : boolean;
  signal SUB_u16_u16_1153_inst_ack_0 : boolean;
  signal SUB_u16_u16_1153_inst_req_1 : boolean;
  signal SUB_u16_u16_1153_inst_ack_1 : boolean;
  signal type_cast_1408_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1436_inst_ack_0 : boolean;
  signal do_while_stmt_956_branch_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1436_inst_req_0 : boolean;
  signal do_while_stmt_956_branch_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1 : boolean;
  signal call_stmt_1170_call_req_0 : boolean;
  signal call_stmt_1170_call_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_req_1 : boolean;
  signal type_cast_887_inst_ack_0 : boolean;
  signal call_stmt_1170_call_req_1 : boolean;
  signal call_stmt_1170_call_ack_1 : boolean;
  signal type_cast_887_inst_req_0 : boolean;
  signal type_cast_1175_inst_req_0 : boolean;
  signal type_cast_1175_inst_ack_0 : boolean;
  signal type_cast_1175_inst_req_1 : boolean;
  signal type_cast_1175_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1433_inst_ack_1 : boolean;
  signal type_cast_1180_inst_req_0 : boolean;
  signal type_cast_1180_inst_ack_0 : boolean;
  signal type_cast_1180_inst_req_1 : boolean;
  signal type_cast_1180_inst_ack_1 : boolean;
  signal phi_stmt_452_ack_0 : boolean;
  signal type_cast_1398_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1433_inst_req_1 : boolean;
  signal type_cast_1190_inst_req_0 : boolean;
  signal type_cast_1190_inst_ack_0 : boolean;
  signal type_cast_1190_inst_req_1 : boolean;
  signal type_cast_1190_inst_ack_1 : boolean;
  signal type_cast_1398_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1433_inst_ack_0 : boolean;
  signal type_cast_1200_inst_req_0 : boolean;
  signal type_cast_1200_inst_ack_0 : boolean;
  signal type_cast_1200_inst_req_1 : boolean;
  signal type_cast_1200_inst_ack_1 : boolean;
  signal phi_stmt_452_req_1 : boolean;
  signal type_cast_1398_inst_ack_0 : boolean;
  signal type_cast_458_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1433_inst_req_0 : boolean;
  signal type_cast_1210_inst_req_0 : boolean;
  signal type_cast_1210_inst_ack_0 : boolean;
  signal type_cast_1210_inst_req_1 : boolean;
  signal if_stmt_1465_branch_ack_0 : boolean;
  signal type_cast_1210_inst_ack_1 : boolean;
  signal type_cast_1398_inst_req_0 : boolean;
  signal type_cast_458_inst_req_1 : boolean;
  signal type_cast_1220_inst_req_0 : boolean;
  signal type_cast_1220_inst_ack_0 : boolean;
  signal type_cast_1220_inst_req_1 : boolean;
  signal type_cast_1220_inst_ack_1 : boolean;
  signal type_cast_458_inst_ack_0 : boolean;
  signal type_cast_1230_inst_req_0 : boolean;
  signal type_cast_1230_inst_ack_0 : boolean;
  signal type_cast_1230_inst_req_1 : boolean;
  signal type_cast_1230_inst_ack_1 : boolean;
  signal type_cast_1240_inst_req_0 : boolean;
  signal type_cast_1240_inst_ack_0 : boolean;
  signal type_cast_1240_inst_req_1 : boolean;
  signal type_cast_1240_inst_ack_1 : boolean;
  signal type_cast_1250_inst_req_0 : boolean;
  signal type_cast_1250_inst_ack_0 : boolean;
  signal type_cast_1250_inst_req_1 : boolean;
  signal type_cast_1250_inst_ack_1 : boolean;
  signal type_cast_1260_inst_req_0 : boolean;
  signal type_cast_1260_inst_ack_0 : boolean;
  signal type_cast_1260_inst_req_1 : boolean;
  signal type_cast_1260_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1262_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1262_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1262_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1262_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1265_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1265_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1265_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1265_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1268_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1268_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1268_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1268_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1271_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1271_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1271_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1271_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1274_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1274_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1274_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1274_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1277_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1277_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1277_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1277_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_ack_1 : boolean;
  signal if_stmt_1293_branch_req_0 : boolean;
  signal if_stmt_1293_branch_ack_1 : boolean;
  signal if_stmt_1293_branch_ack_0 : boolean;
  signal type_cast_1320_inst_req_0 : boolean;
  signal type_cast_1320_inst_ack_0 : boolean;
  signal type_cast_1320_inst_req_1 : boolean;
  signal type_cast_1320_inst_ack_1 : boolean;
  signal array_obj_ref_1349_index_offset_req_0 : boolean;
  signal array_obj_ref_1349_index_offset_ack_0 : boolean;
  signal array_obj_ref_1349_index_offset_req_1 : boolean;
  signal array_obj_ref_1349_index_offset_ack_1 : boolean;
  signal addr_of_1350_final_reg_req_0 : boolean;
  signal addr_of_1350_final_reg_ack_0 : boolean;
  signal addr_of_1350_final_reg_req_1 : boolean;
  signal addr_of_1350_final_reg_ack_1 : boolean;
  signal ptr_deref_1354_load_0_req_0 : boolean;
  signal ptr_deref_1354_load_0_ack_0 : boolean;
  signal ptr_deref_1354_load_0_req_1 : boolean;
  signal ptr_deref_1354_load_0_ack_1 : boolean;
  signal type_cast_1358_inst_req_0 : boolean;
  signal type_cast_1358_inst_ack_0 : boolean;
  signal type_cast_1358_inst_req_1 : boolean;
  signal type_cast_1358_inst_ack_1 : boolean;
  signal phi_stmt_1337_req_0 : boolean;
  signal type_cast_1343_inst_req_0 : boolean;
  signal type_cast_1343_inst_ack_0 : boolean;
  signal type_cast_1343_inst_req_1 : boolean;
  signal type_cast_1343_inst_ack_1 : boolean;
  signal phi_stmt_1337_req_1 : boolean;
  signal phi_stmt_1337_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "ct_core_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  ct_core_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "ct_core_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ct_core_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= ct_core_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ct_core_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  ct_core_CP_34: Block -- control-path 
    signal ct_core_CP_34_elements: BooleanArray(522 downto 0);
    -- 
  begin -- 
    ct_core_CP_34_elements(0) <= ct_core_CP_34_start;
    ct_core_CP_34_symbol <= ct_core_CP_34_elements(522);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	53 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	100 
    -- CP-element group 0: 	103 
    -- CP-element group 0: 	106 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	112 
    -- CP-element group 0: 	115 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	33 
    -- CP-element group 0:  members (98) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_25/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/branch_block_stmt_25__entry__
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392__entry__
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_update_start_
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_Update/cr
      -- 
    cr_183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_45_inst_req_1); -- 
    rr_136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => RPIPE_ConvTranspose_input_pipe_27_inst_req_0); -- 
    cr_155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_32_inst_req_1); -- 
    cr_211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_57_inst_req_1); -- 
    cr_239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_70_inst_req_1); -- 
    cr_267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_82_inst_req_1); -- 
    cr_295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_95_inst_req_1); -- 
    cr_323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_107_inst_req_1); -- 
    cr_351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_120_inst_req_1); -- 
    cr_379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_132_inst_req_1); -- 
    cr_799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_320_inst_req_1); -- 
    cr_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_145_inst_req_1); -- 
    cr_435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_157_inst_req_1); -- 
    cr_463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_170_inst_req_1); -- 
    cr_491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_182_inst_req_1); -- 
    cr_519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_195_inst_req_1); -- 
    cr_547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_207_inst_req_1); -- 
    cr_575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_220_inst_req_1); -- 
    cr_603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_232_inst_req_1); -- 
    cr_631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_245_inst_req_1); -- 
    cr_659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_257_inst_req_1); -- 
    cr_687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_270_inst_req_1); -- 
    cr_715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_282_inst_req_1); -- 
    cr_743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_295_inst_req_1); -- 
    cr_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_307_inst_req_1); -- 
    cr_813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_330_inst_req_1); -- 
    cr_827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_339_inst_req_1); -- 
    cr_841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_358_inst_req_1); -- 
    cr_855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_362_inst_req_1); -- 
    cr_869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_371_inst_req_1); -- 
    cr_883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(0), ack => type_cast_380_inst_req_1); -- 
    -- CP-element group 1:  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	396 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	400 
    -- CP-element group 1: 	402 
    -- CP-element group 1: 	397 
    -- CP-element group 1: 	398 
    -- CP-element group 1: 	399 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_25/do_while_stmt_956__exit__
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186__entry__
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/$entry
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_update_start_
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_Sample/crr
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_Update/ccr
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_update_start_
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_update_start_
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_Update/cr
      -- 
    crr_2407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(1), ack => call_stmt_1170_call_req_0); -- 
    ccr_2412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(1), ack => call_stmt_1170_call_req_1); -- 
    rr_2421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(1), ack => type_cast_1175_inst_req_0); -- 
    cr_2426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(1), ack => type_cast_1175_inst_req_1); -- 
    cr_2440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(1), ack => type_cast_1180_inst_req_1); -- 
    ct_core_CP_34_elements(1) <= ct_core_CP_34_elements(396);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_update_start_
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_Update/cr
      -- 
    ra_137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_27_inst_ack_0, ack => ct_core_CP_34_elements(2)); -- 
    cr_141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(2), ack => RPIPE_ConvTranspose_input_pipe_27_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_27_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_Sample/rr
      -- 
    ca_142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_27_inst_ack_1, ack => ct_core_CP_34_elements(3)); -- 
    rr_150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(3), ack => type_cast_32_inst_req_0); -- 
    rr_164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(3), ack => RPIPE_ConvTranspose_input_pipe_41_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_Sample/ra
      -- 
    ra_151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_32_inst_ack_0, ack => ct_core_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	101 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_32_Update/ca
      -- 
    ca_156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_32_inst_ack_1, ack => ct_core_CP_34_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_update_start_
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_Update/cr
      -- 
    ra_165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_41_inst_ack_0, ack => ct_core_CP_34_elements(6)); -- 
    cr_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(6), ack => RPIPE_ConvTranspose_input_pipe_41_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_41_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_Sample/rr
      -- 
    ca_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_41_inst_ack_1, ack => ct_core_CP_34_elements(7)); -- 
    rr_178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(7), ack => type_cast_45_inst_req_0); -- 
    rr_192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(7), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_Sample/$exit
      -- 
    ra_179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_45_inst_ack_0, ack => ct_core_CP_34_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	101 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_45_update_completed_
      -- 
    ca_184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_45_inst_ack_1, ack => ct_core_CP_34_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_update_start_
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_Update/cr
      -- 
    ra_193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_0, ack => ct_core_CP_34_elements(10)); -- 
    cr_197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(10), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_53_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_Sample/rr
      -- 
    ca_198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_1, ack => ct_core_CP_34_elements(11)); -- 
    rr_206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(11), ack => type_cast_57_inst_req_0); -- 
    rr_220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(11), ack => RPIPE_ConvTranspose_input_pipe_66_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_Sample/ra
      -- 
    ra_207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_0, ack => ct_core_CP_34_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	101 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_57_Update/ca
      -- 
    ca_212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_1, ack => ct_core_CP_34_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_update_start_
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_Update/cr
      -- 
    ra_221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_66_inst_ack_0, ack => ct_core_CP_34_elements(14)); -- 
    cr_225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(14), ack => RPIPE_ConvTranspose_input_pipe_66_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_66_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_Sample/rr
      -- 
    ca_226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_66_inst_ack_1, ack => ct_core_CP_34_elements(15)); -- 
    rr_234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(15), ack => type_cast_70_inst_req_0); -- 
    rr_248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(15), ack => RPIPE_ConvTranspose_input_pipe_78_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_Sample/ra
      -- 
    ra_235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_70_inst_ack_0, ack => ct_core_CP_34_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	101 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_70_Update/ca
      -- 
    ca_240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_70_inst_ack_1, ack => ct_core_CP_34_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_update_start_
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_Update/cr
      -- 
    ra_249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_78_inst_ack_0, ack => ct_core_CP_34_elements(18)); -- 
    cr_253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(18), ack => RPIPE_ConvTranspose_input_pipe_78_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_78_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_Sample/rr
      -- 
    ca_254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_78_inst_ack_1, ack => ct_core_CP_34_elements(19)); -- 
    rr_262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(19), ack => type_cast_82_inst_req_0); -- 
    rr_276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(19), ack => RPIPE_ConvTranspose_input_pipe_91_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_Sample/ra
      -- 
    ra_263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_0, ack => ct_core_CP_34_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	98 
    -- CP-element group 21: 	110 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_82_Update/ca
      -- 
    ca_268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_1, ack => ct_core_CP_34_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_update_start_
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_Update/cr
      -- 
    ra_277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_91_inst_ack_0, ack => ct_core_CP_34_elements(22)); -- 
    cr_281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(22), ack => RPIPE_ConvTranspose_input_pipe_91_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_91_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_Sample/rr
      -- 
    ca_282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_91_inst_ack_1, ack => ct_core_CP_34_elements(23)); -- 
    rr_290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(23), ack => type_cast_95_inst_req_0); -- 
    rr_304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(23), ack => RPIPE_ConvTranspose_input_pipe_103_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_Sample/ra
      -- 
    ra_291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_0, ack => ct_core_CP_34_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	98 
    -- CP-element group 25: 	110 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_95_Update/ca
      -- 
    ca_296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_1, ack => ct_core_CP_34_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_update_start_
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_Update/cr
      -- 
    ra_305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_103_inst_ack_0, ack => ct_core_CP_34_elements(26)); -- 
    cr_309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(26), ack => RPIPE_ConvTranspose_input_pipe_103_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_103_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_Sample/rr
      -- 
    ca_310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_103_inst_ack_1, ack => ct_core_CP_34_elements(27)); -- 
    rr_318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(27), ack => type_cast_107_inst_req_0); -- 
    rr_332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(27), ack => RPIPE_ConvTranspose_input_pipe_116_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_Sample/ra
      -- 
    ra_319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_0, ack => ct_core_CP_34_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	104 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_107_Update/ca
      -- 
    ca_324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_1, ack => ct_core_CP_34_elements(29)); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_update_start_
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_Update/cr
      -- 
    ra_333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_116_inst_ack_0, ack => ct_core_CP_34_elements(30)); -- 
    cr_337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(30), ack => RPIPE_ConvTranspose_input_pipe_116_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_116_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_Sample/rr
      -- 
    ca_338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_116_inst_ack_1, ack => ct_core_CP_34_elements(31)); -- 
    rr_346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(31), ack => type_cast_120_inst_req_0); -- 
    rr_360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(31), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_Sample/ra
      -- 
    ra_347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_0, ack => ct_core_CP_34_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	104 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_120_Update/ca
      -- 
    ca_352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_120_inst_ack_1, ack => ct_core_CP_34_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_update_start_
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_Update/cr
      -- 
    ra_361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_0, ack => ct_core_CP_34_elements(34)); -- 
    cr_365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(34), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_128_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_Sample/rr
      -- 
    ca_366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_1, ack => ct_core_CP_34_elements(35)); -- 
    rr_388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(35), ack => RPIPE_ConvTranspose_input_pipe_141_inst_req_0); -- 
    rr_374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(35), ack => type_cast_132_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_Sample/ra
      -- 
    ra_375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_132_inst_ack_0, ack => ct_core_CP_34_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	104 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_132_Update/ca
      -- 
    ca_380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_132_inst_ack_1, ack => ct_core_CP_34_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_update_start_
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_Update/cr
      -- 
    ra_389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_141_inst_ack_0, ack => ct_core_CP_34_elements(38)); -- 
    cr_393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(38), ack => RPIPE_ConvTranspose_input_pipe_141_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_141_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_Sample/rr
      -- 
    ca_394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_141_inst_ack_1, ack => ct_core_CP_34_elements(39)); -- 
    rr_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(39), ack => type_cast_145_inst_req_0); -- 
    rr_416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(39), ack => RPIPE_ConvTranspose_input_pipe_153_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_Sample/ra
      -- 
    ra_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_0, ack => ct_core_CP_34_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	104 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_145_Update/ca
      -- 
    ca_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_145_inst_ack_1, ack => ct_core_CP_34_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_update_start_
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_Update/cr
      -- 
    ra_417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_153_inst_ack_0, ack => ct_core_CP_34_elements(42)); -- 
    cr_421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(42), ack => RPIPE_ConvTranspose_input_pipe_153_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_153_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_Sample/rr
      -- 
    ca_422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_153_inst_ack_1, ack => ct_core_CP_34_elements(43)); -- 
    rr_430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(43), ack => type_cast_157_inst_req_0); -- 
    rr_444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(43), ack => RPIPE_ConvTranspose_input_pipe_166_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_Sample/ra
      -- 
    ra_431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_0, ack => ct_core_CP_34_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	107 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_157_Update/ca
      -- 
    ca_436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_1, ack => ct_core_CP_34_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_update_start_
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_Update/cr
      -- 
    ra_445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_166_inst_ack_0, ack => ct_core_CP_34_elements(46)); -- 
    cr_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(46), ack => RPIPE_ConvTranspose_input_pipe_166_inst_req_1); -- 
    -- CP-element group 47:  fork  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	50 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_166_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_Sample/rr
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_Sample/rr
      -- 
    ca_450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_166_inst_ack_1, ack => ct_core_CP_34_elements(47)); -- 
    rr_472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(47), ack => RPIPE_ConvTranspose_input_pipe_178_inst_req_0); -- 
    rr_458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(47), ack => type_cast_170_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_Sample/ra
      -- 
    ra_459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_170_inst_ack_0, ack => ct_core_CP_34_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	107 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_170_Update/ca
      -- 
    ca_464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_170_inst_ack_1, ack => ct_core_CP_34_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	47 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_update_start_
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_Update/cr
      -- 
    ra_473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_178_inst_ack_0, ack => ct_core_CP_34_elements(50)); -- 
    cr_477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(50), ack => RPIPE_ConvTranspose_input_pipe_178_inst_req_1); -- 
    -- CP-element group 51:  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_178_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_Sample/rr
      -- 
    ca_478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_178_inst_ack_1, ack => ct_core_CP_34_elements(51)); -- 
    rr_500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(51), ack => RPIPE_ConvTranspose_input_pipe_191_inst_req_0); -- 
    rr_486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(51), ack => type_cast_182_inst_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_Sample/ra
      -- 
    ra_487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_0, ack => ct_core_CP_34_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	0 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	107 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_182_Update/ca
      -- 
    ca_492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_1, ack => ct_core_CP_34_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_update_start_
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_Update/cr
      -- 
    ra_501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_191_inst_ack_0, ack => ct_core_CP_34_elements(54)); -- 
    cr_505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(54), ack => RPIPE_ConvTranspose_input_pipe_191_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_191_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_Sample/rr
      -- 
    ca_506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_191_inst_ack_1, ack => ct_core_CP_34_elements(55)); -- 
    rr_514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(55), ack => type_cast_195_inst_req_0); -- 
    rr_528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(55), ack => RPIPE_ConvTranspose_input_pipe_203_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_Sample/ra
      -- 
    ra_515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_195_inst_ack_0, ack => ct_core_CP_34_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	107 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_195_Update/ca
      -- 
    ca_520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_195_inst_ack_1, ack => ct_core_CP_34_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_update_start_
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_Update/cr
      -- 
    ra_529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_203_inst_ack_0, ack => ct_core_CP_34_elements(58)); -- 
    cr_533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(58), ack => RPIPE_ConvTranspose_input_pipe_203_inst_req_1); -- 
    -- CP-element group 59:  fork  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	62 
    -- CP-element group 59:  members (9) 
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_203_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_Sample/rr
      -- 
    ca_534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_203_inst_ack_1, ack => ct_core_CP_34_elements(59)); -- 
    rr_542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(59), ack => type_cast_207_inst_req_0); -- 
    rr_556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(59), ack => RPIPE_ConvTranspose_input_pipe_216_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_Sample/ra
      -- 
    ra_543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_207_inst_ack_0, ack => ct_core_CP_34_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	116 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_207_Update/ca
      -- 
    ca_548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_207_inst_ack_1, ack => ct_core_CP_34_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_update_start_
      -- CP-element group 62: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_Update/cr
      -- 
    ra_557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_216_inst_ack_0, ack => ct_core_CP_34_elements(62)); -- 
    cr_561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(62), ack => RPIPE_ConvTranspose_input_pipe_216_inst_req_1); -- 
    -- CP-element group 63:  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_216_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_Sample/rr
      -- 
    ca_562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_216_inst_ack_1, ack => ct_core_CP_34_elements(63)); -- 
    rr_570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(63), ack => type_cast_220_inst_req_0); -- 
    rr_584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(63), ack => RPIPE_ConvTranspose_input_pipe_228_inst_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_Sample/ra
      -- 
    ra_571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_0, ack => ct_core_CP_34_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	116 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_220_Update/ca
      -- 
    ca_576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_1, ack => ct_core_CP_34_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_update_start_
      -- CP-element group 66: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_Update/cr
      -- 
    ra_585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_228_inst_ack_0, ack => ct_core_CP_34_elements(66)); -- 
    cr_589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(66), ack => RPIPE_ConvTranspose_input_pipe_228_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	70 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_228_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_Sample/rr
      -- 
    ca_590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_228_inst_ack_1, ack => ct_core_CP_34_elements(67)); -- 
    rr_598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(67), ack => type_cast_232_inst_req_0); -- 
    rr_612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(67), ack => RPIPE_ConvTranspose_input_pipe_241_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_Sample/ra
      -- 
    ra_599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_232_inst_ack_0, ack => ct_core_CP_34_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	116 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_232_Update/ca
      -- 
    ca_604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_232_inst_ack_1, ack => ct_core_CP_34_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_update_start_
      -- CP-element group 70: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_Update/cr
      -- 
    ra_613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_241_inst_ack_0, ack => ct_core_CP_34_elements(70)); -- 
    cr_617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(70), ack => RPIPE_ConvTranspose_input_pipe_241_inst_req_1); -- 
    -- CP-element group 71:  fork  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	74 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_241_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_Sample/rr
      -- 
    ca_618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_241_inst_ack_1, ack => ct_core_CP_34_elements(71)); -- 
    rr_626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(71), ack => type_cast_245_inst_req_0); -- 
    rr_640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(71), ack => RPIPE_ConvTranspose_input_pipe_253_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_Sample/ra
      -- 
    ra_627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_245_inst_ack_0, ack => ct_core_CP_34_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	116 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_245_Update/ca
      -- 
    ca_632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_245_inst_ack_1, ack => ct_core_CP_34_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	71 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_update_start_
      -- CP-element group 74: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_Update/cr
      -- 
    ra_641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_253_inst_ack_0, ack => ct_core_CP_34_elements(74)); -- 
    cr_645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(74), ack => RPIPE_ConvTranspose_input_pipe_253_inst_req_1); -- 
    -- CP-element group 75:  fork  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (9) 
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_253_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_Sample/rr
      -- 
    ca_646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_253_inst_ack_1, ack => ct_core_CP_34_elements(75)); -- 
    rr_668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(75), ack => RPIPE_ConvTranspose_input_pipe_266_inst_req_0); -- 
    rr_654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(75), ack => type_cast_257_inst_req_0); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_Sample/ra
      -- 
    ra_655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_257_inst_ack_0, ack => ct_core_CP_34_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	113 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_257_Update/ca
      -- 
    ca_660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_257_inst_ack_1, ack => ct_core_CP_34_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_update_start_
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_Update/cr
      -- 
    ra_669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_266_inst_ack_0, ack => ct_core_CP_34_elements(78)); -- 
    cr_673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(78), ack => RPIPE_ConvTranspose_input_pipe_266_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_266_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_Sample/rr
      -- 
    ca_674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_266_inst_ack_1, ack => ct_core_CP_34_elements(79)); -- 
    rr_682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(79), ack => type_cast_270_inst_req_0); -- 
    rr_696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(79), ack => RPIPE_ConvTranspose_input_pipe_278_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_Sample/ra
      -- 
    ra_683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_270_inst_ack_0, ack => ct_core_CP_34_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	113 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_270_Update/ca
      -- 
    ca_688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_270_inst_ack_1, ack => ct_core_CP_34_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_update_start_
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_Update/cr
      -- 
    ra_697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_278_inst_ack_0, ack => ct_core_CP_34_elements(82)); -- 
    cr_701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(82), ack => RPIPE_ConvTranspose_input_pipe_278_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_278_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_Sample/rr
      -- 
    ca_702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_278_inst_ack_1, ack => ct_core_CP_34_elements(83)); -- 
    rr_710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(83), ack => type_cast_282_inst_req_0); -- 
    rr_724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(83), ack => RPIPE_ConvTranspose_input_pipe_291_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_Sample/ra
      -- 
    ra_711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_282_inst_ack_0, ack => ct_core_CP_34_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	113 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_282_Update/ca
      -- 
    ca_716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_282_inst_ack_1, ack => ct_core_CP_34_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_update_start_
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_Update/cr
      -- 
    ra_725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_291_inst_ack_0, ack => ct_core_CP_34_elements(86)); -- 
    cr_729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(86), ack => RPIPE_ConvTranspose_input_pipe_291_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_291_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_Sample/rr
      -- 
    ca_730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_291_inst_ack_1, ack => ct_core_CP_34_elements(87)); -- 
    rr_738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(87), ack => type_cast_295_inst_req_0); -- 
    rr_752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(87), ack => RPIPE_ConvTranspose_input_pipe_303_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_Sample/ra
      -- 
    ra_739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_295_inst_ack_0, ack => ct_core_CP_34_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	113 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_295_Update/ca
      -- 
    ca_744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_295_inst_ack_1, ack => ct_core_CP_34_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_update_start_
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_Update/cr
      -- 
    ra_753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_303_inst_ack_0, ack => ct_core_CP_34_elements(90)); -- 
    cr_757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(90), ack => RPIPE_ConvTranspose_input_pipe_303_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_303_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_Sample/$entry
      -- 
    ca_758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_303_inst_ack_1, ack => ct_core_CP_34_elements(91)); -- 
    rr_766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(91), ack => type_cast_307_inst_req_0); -- 
    rr_780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(91), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_Sample/ra
      -- 
    ra_767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_307_inst_ack_0, ack => ct_core_CP_34_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	116 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_307_Update/ca
      -- 
    ca_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_307_inst_ack_1, ack => ct_core_CP_34_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_update_start_
      -- CP-element group 94: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_Sample/$exit
      -- 
    ra_781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_0, ack => ct_core_CP_34_elements(94)); -- 
    cr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(94), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_1); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/RPIPE_ConvTranspose_input_pipe_316_update_completed_
      -- 
    ca_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_1, ack => ct_core_CP_34_elements(95)); -- 
    rr_794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(95), ack => type_cast_320_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_Sample/ra
      -- 
    ra_795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_0, ack => ct_core_CP_34_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	116 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_320_Update/ca
      -- 
    ca_800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_1, ack => ct_core_CP_34_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	21 
    -- CP-element group 98: 	25 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_Sample/rr
      -- 
    rr_808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(98), ack => type_cast_330_inst_req_0); -- 
    ct_core_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "ct_core_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(21) & ct_core_CP_34_elements(25);
      gj_ct_core_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_Sample/ra
      -- 
    ra_809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_330_inst_ack_0, ack => ct_core_CP_34_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	0 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	116 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_330_Update/ca
      -- 
    ca_814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_330_inst_ack_1, ack => ct_core_CP_34_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	5 
    -- CP-element group 101: 	9 
    -- CP-element group 101: 	13 
    -- CP-element group 101: 	17 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_Sample/rr
      -- 
    rr_822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(101), ack => type_cast_339_inst_req_0); -- 
    ct_core_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(5) & ct_core_CP_34_elements(9) & ct_core_CP_34_elements(13) & ct_core_CP_34_elements(17);
      gj_ct_core_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_Sample/ra
      -- 
    ra_823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_339_inst_ack_0, ack => ct_core_CP_34_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	0 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	116 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_339_Update/ca
      -- 
    ca_828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_339_inst_ack_1, ack => ct_core_CP_34_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	41 
    -- CP-element group 104: 	37 
    -- CP-element group 104: 	29 
    -- CP-element group 104: 	33 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_Sample/rr
      -- 
    rr_836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(104), ack => type_cast_358_inst_req_0); -- 
    ct_core_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(41) & ct_core_CP_34_elements(37) & ct_core_CP_34_elements(29) & ct_core_CP_34_elements(33);
      gj_ct_core_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_Sample/ra
      -- 
    ra_837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_0, ack => ct_core_CP_34_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	0 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	116 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_358_Update/ca
      -- 
    ca_842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_1, ack => ct_core_CP_34_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	57 
    -- CP-element group 107: 	53 
    -- CP-element group 107: 	45 
    -- CP-element group 107: 	49 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_Sample/rr
      -- 
    rr_850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(107), ack => type_cast_362_inst_req_0); -- 
    ct_core_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(57) & ct_core_CP_34_elements(53) & ct_core_CP_34_elements(45) & ct_core_CP_34_elements(49);
      gj_ct_core_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_Sample/ra
      -- 
    ra_851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_362_inst_ack_0, ack => ct_core_CP_34_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	116 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_362_Update/ca
      -- 
    ca_856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_362_inst_ack_1, ack => ct_core_CP_34_elements(109)); -- 
    -- CP-element group 110:  join  transition  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	21 
    -- CP-element group 110: 	25 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_Sample/rr
      -- 
    rr_864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(110), ack => type_cast_371_inst_req_0); -- 
    ct_core_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(21) & ct_core_CP_34_elements(25);
      gj_ct_core_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_Sample/ra
      -- 
    ra_865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_0, ack => ct_core_CP_34_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	0 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	116 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_371_Update/ca
      -- 
    ca_870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_1, ack => ct_core_CP_34_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	77 
    -- CP-element group 113: 	85 
    -- CP-element group 113: 	89 
    -- CP-element group 113: 	81 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_Sample/rr
      -- 
    rr_878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(113), ack => type_cast_380_inst_req_0); -- 
    ct_core_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(77) & ct_core_CP_34_elements(85) & ct_core_CP_34_elements(89) & ct_core_CP_34_elements(81);
      gj_ct_core_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_Sample/ra
      -- 
    ra_879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_0, ack => ct_core_CP_34_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	0 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/type_cast_380_Update/ca
      -- 
    ca_884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_380_inst_ack_1, ack => ct_core_CP_34_elements(115)); -- 
    -- CP-element group 116:  branch  join  transition  place  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	61 
    -- CP-element group 116: 	65 
    -- CP-element group 116: 	69 
    -- CP-element group 116: 	73 
    -- CP-element group 116: 	93 
    -- CP-element group 116: 	97 
    -- CP-element group 116: 	100 
    -- CP-element group 116: 	103 
    -- CP-element group 116: 	106 
    -- CP-element group 116: 	109 
    -- CP-element group 116: 	112 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (10) 
      -- CP-element group 116: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392__exit__
      -- CP-element group 116: 	 branch_block_stmt_25/if_stmt_393__entry__
      -- CP-element group 116: 	 branch_block_stmt_25/assign_stmt_28_to_assign_stmt_392/$exit
      -- CP-element group 116: 	 branch_block_stmt_25/if_stmt_393_dead_link/$entry
      -- CP-element group 116: 	 branch_block_stmt_25/if_stmt_393_eval_test/$entry
      -- CP-element group 116: 	 branch_block_stmt_25/if_stmt_393_eval_test/$exit
      -- CP-element group 116: 	 branch_block_stmt_25/if_stmt_393_eval_test/branch_req
      -- CP-element group 116: 	 branch_block_stmt_25/R_cmp467_394_place
      -- CP-element group 116: 	 branch_block_stmt_25/if_stmt_393_if_link/$entry
      -- CP-element group 116: 	 branch_block_stmt_25/if_stmt_393_else_link/$entry
      -- 
    branch_req_892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(116), ack => if_stmt_393_branch_req_0); -- 
    ct_core_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(61) & ct_core_CP_34_elements(65) & ct_core_CP_34_elements(69) & ct_core_CP_34_elements(73) & ct_core_CP_34_elements(93) & ct_core_CP_34_elements(97) & ct_core_CP_34_elements(100) & ct_core_CP_34_elements(103) & ct_core_CP_34_elements(106) & ct_core_CP_34_elements(109) & ct_core_CP_34_elements(112) & ct_core_CP_34_elements(115);
      gj_ct_core_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	121 
    -- CP-element group 117: 	122 
    -- CP-element group 117:  members (18) 
      -- CP-element group 117: 	 branch_block_stmt_25/merge_stmt_414__exit__
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449__entry__
      -- CP-element group 117: 	 branch_block_stmt_25/if_stmt_393_if_link/$exit
      -- CP-element group 117: 	 branch_block_stmt_25/if_stmt_393_if_link/if_choice_transition
      -- CP-element group 117: 	 branch_block_stmt_25/entry_bbx_xnph469
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/$entry
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_update_start_
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_Update/cr
      -- CP-element group 117: 	 branch_block_stmt_25/merge_stmt_414_PhiAck/dummy
      -- CP-element group 117: 	 branch_block_stmt_25/merge_stmt_414_PhiAck/$exit
      -- CP-element group 117: 	 branch_block_stmt_25/merge_stmt_414_PhiAck/$entry
      -- CP-element group 117: 	 branch_block_stmt_25/entry_bbx_xnph469_PhiReq/$exit
      -- CP-element group 117: 	 branch_block_stmt_25/entry_bbx_xnph469_PhiReq/$entry
      -- CP-element group 117: 	 branch_block_stmt_25/merge_stmt_414_PhiReqMerge
      -- 
    if_choice_transition_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_393_branch_ack_1, ack => ct_core_CP_34_elements(117)); -- 
    rr_936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(117), ack => type_cast_435_inst_req_0); -- 
    cr_941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(117), ack => type_cast_435_inst_req_1); -- 
    -- CP-element group 118:  transition  place  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	495 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_25/if_stmt_393_else_link/$exit
      -- CP-element group 118: 	 branch_block_stmt_25/if_stmt_393_else_link/else_choice_transition
      -- CP-element group 118: 	 branch_block_stmt_25/entry_forx_xcond171x_xpreheader
      -- CP-element group 118: 	 branch_block_stmt_25/entry_forx_xcond171x_xpreheader_PhiReq/$exit
      -- CP-element group 118: 	 branch_block_stmt_25/entry_forx_xcond171x_xpreheader_PhiReq/$entry
      -- 
    else_choice_transition_901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_393_branch_ack_0, ack => ct_core_CP_34_elements(118)); -- 
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	495 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	165 
    -- CP-element group 119: 	166 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_25/merge_stmt_621__exit__
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656__entry__
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_update_start_
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/$entry
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_25/if_stmt_408_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_25/if_stmt_408_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_25/forx_xcond171x_xpreheader_bbx_xnph465
      -- CP-element group 119: 	 branch_block_stmt_25/merge_stmt_621_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_25/merge_stmt_621_PhiAck/dummy
      -- CP-element group 119: 	 branch_block_stmt_25/merge_stmt_621_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_25/merge_stmt_621_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_25/forx_xcond171x_xpreheader_bbx_xnph465_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_25/forx_xcond171x_xpreheader_bbx_xnph465_PhiReq/$entry
      -- 
    if_choice_transition_919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_408_branch_ack_1, ack => ct_core_CP_34_elements(119)); -- 
    rr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(119), ack => type_cast_642_inst_req_0); -- 
    cr_1300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(119), ack => type_cast_642_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	495 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	508 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_25/forx_xcond171x_xpreheader_forx_xend231_PhiReq/$exit
      -- CP-element group 120: 	 branch_block_stmt_25/if_stmt_408_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_25/if_stmt_408_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_25/forx_xcond171x_xpreheader_forx_xend231
      -- CP-element group 120: 	 branch_block_stmt_25/forx_xcond171x_xpreheader_forx_xend231_PhiReq/$entry
      -- 
    else_choice_transition_923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_408_branch_ack_0, ack => ct_core_CP_34_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	117 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_Sample/ra
      -- 
    ra_937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_435_inst_ack_0, ack => ct_core_CP_34_elements(121)); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	117 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	496 
    -- CP-element group 122:  members (9) 
      -- CP-element group 122: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449__exit__
      -- CP-element group 122: 	 branch_block_stmt_25/bbx_xnph469_forx_xbody
      -- CP-element group 122: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/$exit
      -- CP-element group 122: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_25/assign_stmt_420_to_assign_stmt_449/type_cast_435_Update/ca
      -- CP-element group 122: 	 branch_block_stmt_25/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/$entry
      -- CP-element group 122: 	 branch_block_stmt_25/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_452/$entry
      -- CP-element group 122: 	 branch_block_stmt_25/bbx_xnph469_forx_xbody_PhiReq/$entry
      -- 
    ca_942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_435_inst_ack_1, ack => ct_core_CP_34_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	501 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	162 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_final_index_sum_regn_Sample/ack
      -- CP-element group 123: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_final_index_sum_regn_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_final_index_sum_regn_sample_complete
      -- 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_464_index_offset_ack_0, ack => ct_core_CP_34_elements(123)); -- 
    -- CP-element group 124:  transition  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	501 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (11) 
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_base_plus_offset/sum_rename_req
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_base_plus_offset/$exit
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_base_plus_offset/$entry
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_final_index_sum_regn_Update/ack
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_final_index_sum_regn_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_request/req
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_request/$entry
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_base_plus_offset/sum_rename_ack
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_root_address_calculated
      -- CP-element group 124: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_offset_calculated
      -- 
    ack_976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_464_index_offset_ack_1, ack => ct_core_CP_34_elements(124)); -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(124), ack => addr_of_465_final_reg_req_0); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_request/ack
      -- CP-element group 125: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_request/$exit
      -- CP-element group 125: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_sample_completed_
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_465_final_reg_ack_0, ack => ct_core_CP_34_elements(125)); -- 
    -- CP-element group 126:  fork  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	501 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	159 
    -- CP-element group 126:  members (19) 
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_word_addrgen/root_register_req
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_word_addrgen/$exit
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_word_addrgen/$entry
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_base_addr_resize/base_resize_ack
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_base_addr_resize/base_resize_req
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_base_addr_resize/$exit
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_base_addr_resize/$entry
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_base_address_resized
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_word_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_base_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_word_addrgen/root_register_ack
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_complete/ack
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_complete/$exit
      -- CP-element group 126: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_update_completed_
      -- 
    ack_991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_465_final_reg_ack_1, ack => ct_core_CP_34_elements(126)); -- 
    -- CP-element group 127:  transition  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	501 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (6) 
      -- CP-element group 127: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_update_start_
      -- CP-element group 127: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_Update/cr
      -- CP-element group 127: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_Sample/ra
      -- CP-element group 127: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_sample_completed_
      -- 
    ra_1000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_468_inst_ack_0, ack => ct_core_CP_34_elements(127)); -- 
    cr_1004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(127), ack => RPIPE_ConvTranspose_input_pipe_468_inst_req_1); -- 
    -- CP-element group 128:  fork  transition  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128: 	131 
    -- CP-element group 128:  members (9) 
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_Update/ca
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_update_completed_
      -- 
    ca_1005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_468_inst_ack_1, ack => ct_core_CP_34_elements(128)); -- 
    rr_1013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(128), ack => type_cast_472_inst_req_0); -- 
    rr_1027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(128), ack => RPIPE_ConvTranspose_input_pipe_481_inst_req_0); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_sample_completed_
      -- 
    ra_1014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_472_inst_ack_0, ack => ct_core_CP_34_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	501 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	159 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_update_completed_
      -- 
    ca_1019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_472_inst_ack_1, ack => ct_core_CP_34_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	128 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_update_start_
      -- CP-element group 131: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_sample_completed_
      -- 
    ra_1028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_481_inst_ack_0, ack => ct_core_CP_34_elements(131)); -- 
    cr_1032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(131), ack => RPIPE_ConvTranspose_input_pipe_481_inst_req_1); -- 
    -- CP-element group 132:  fork  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132: 	135 
    -- CP-element group 132:  members (9) 
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_481_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_Sample/rr
      -- 
    ca_1033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_481_inst_ack_1, ack => ct_core_CP_34_elements(132)); -- 
    rr_1041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(132), ack => type_cast_485_inst_req_0); -- 
    rr_1055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(132), ack => RPIPE_ConvTranspose_input_pipe_499_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_Sample/ra
      -- 
    ra_1042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_0, ack => ct_core_CP_34_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	501 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	159 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_Update/$exit
      -- 
    ca_1047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_485_inst_ack_1, ack => ct_core_CP_34_elements(134)); -- 
    -- CP-element group 135:  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	132 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (6) 
      -- CP-element group 135: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_update_start_
      -- CP-element group 135: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_Update/cr
      -- CP-element group 135: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_Sample/ra
      -- 
    ra_1056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_499_inst_ack_0, ack => ct_core_CP_34_elements(135)); -- 
    cr_1060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(135), ack => RPIPE_ConvTranspose_input_pipe_499_inst_req_1); -- 
    -- CP-element group 136:  fork  transition  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136: 	139 
    -- CP-element group 136:  members (9) 
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_Sample/rr
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_Sample/rr
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_499_Update/$exit
      -- 
    ca_1061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_499_inst_ack_1, ack => ct_core_CP_34_elements(136)); -- 
    rr_1069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(136), ack => type_cast_503_inst_req_0); -- 
    rr_1083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(136), ack => RPIPE_ConvTranspose_input_pipe_517_inst_req_0); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_sample_completed_
      -- 
    ra_1070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_503_inst_ack_0, ack => ct_core_CP_34_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	501 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	159 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_update_completed_
      -- 
    ca_1075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_503_inst_ack_1, ack => ct_core_CP_34_elements(138)); -- 
    -- CP-element group 139:  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	136 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139:  members (6) 
      -- CP-element group 139: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_update_start_
      -- CP-element group 139: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_Update/cr
      -- CP-element group 139: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_Sample/ra
      -- 
    ra_1084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_517_inst_ack_0, ack => ct_core_CP_34_elements(139)); -- 
    cr_1088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(139), ack => RPIPE_ConvTranspose_input_pipe_517_inst_req_1); -- 
    -- CP-element group 140:  fork  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140: 	143 
    -- CP-element group 140:  members (9) 
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_Sample/rr
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_Sample/rr
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_517_Update/$exit
      -- 
    ca_1089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_517_inst_ack_1, ack => ct_core_CP_34_elements(140)); -- 
    rr_1097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(140), ack => type_cast_521_inst_req_0); -- 
    rr_1111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(140), ack => RPIPE_ConvTranspose_input_pipe_535_inst_req_0); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_sample_completed_
      -- 
    ra_1098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_521_inst_ack_0, ack => ct_core_CP_34_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	501 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	159 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_update_completed_
      -- 
    ca_1103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_521_inst_ack_1, ack => ct_core_CP_34_elements(142)); -- 
    -- CP-element group 143:  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	140 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (6) 
      -- CP-element group 143: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_Update/cr
      -- CP-element group 143: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_update_start_
      -- CP-element group 143: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_sample_completed_
      -- 
    ra_1112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_535_inst_ack_0, ack => ct_core_CP_34_elements(143)); -- 
    cr_1116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(143), ack => RPIPE_ConvTranspose_input_pipe_535_inst_req_1); -- 
    -- CP-element group 144:  fork  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144: 	147 
    -- CP-element group 144:  members (9) 
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_535_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_sample_start_
      -- 
    ca_1117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_535_inst_ack_1, ack => ct_core_CP_34_elements(144)); -- 
    rr_1125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(144), ack => type_cast_539_inst_req_0); -- 
    rr_1139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(144), ack => RPIPE_ConvTranspose_input_pipe_553_inst_req_0); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_Sample/ra
      -- CP-element group 145: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_sample_completed_
      -- 
    ra_1126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_539_inst_ack_0, ack => ct_core_CP_34_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	501 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	159 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_update_completed_
      -- 
    ca_1131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_539_inst_ack_1, ack => ct_core_CP_34_elements(146)); -- 
    -- CP-element group 147:  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	144 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (6) 
      -- CP-element group 147: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_Update/cr
      -- CP-element group 147: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_update_start_
      -- CP-element group 147: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_sample_completed_
      -- 
    ra_1140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_553_inst_ack_0, ack => ct_core_CP_34_elements(147)); -- 
    cr_1144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(147), ack => RPIPE_ConvTranspose_input_pipe_553_inst_req_1); -- 
    -- CP-element group 148:  fork  transition  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: 	151 
    -- CP-element group 148:  members (9) 
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_Sample/rr
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_Sample/$entry
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_Sample/rr
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_Sample/$entry
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_553_update_completed_
      -- 
    ca_1145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_553_inst_ack_1, ack => ct_core_CP_34_elements(148)); -- 
    rr_1153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(148), ack => type_cast_557_inst_req_0); -- 
    rr_1167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(148), ack => RPIPE_ConvTranspose_input_pipe_571_inst_req_0); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_sample_completed_
      -- 
    ra_1154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_557_inst_ack_0, ack => ct_core_CP_34_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	501 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	159 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_update_completed_
      -- 
    ca_1159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_557_inst_ack_1, ack => ct_core_CP_34_elements(150)); -- 
    -- CP-element group 151:  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	148 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (6) 
      -- CP-element group 151: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_update_start_
      -- CP-element group 151: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_Update/cr
      -- CP-element group 151: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_Update/$entry
      -- 
    ra_1168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_571_inst_ack_0, ack => ct_core_CP_34_elements(151)); -- 
    cr_1172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(151), ack => RPIPE_ConvTranspose_input_pipe_571_inst_req_1); -- 
    -- CP-element group 152:  fork  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152: 	155 
    -- CP-element group 152:  members (9) 
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_Sample/rr
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_Sample/rr
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_571_Update/$exit
      -- 
    ca_1173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_571_inst_ack_1, ack => ct_core_CP_34_elements(152)); -- 
    rr_1181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(152), ack => type_cast_575_inst_req_0); -- 
    rr_1195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(152), ack => RPIPE_ConvTranspose_input_pipe_589_inst_req_0); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_sample_completed_
      -- 
    ra_1182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_575_inst_ack_0, ack => ct_core_CP_34_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	501 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	159 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_update_completed_
      -- 
    ca_1187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_575_inst_ack_1, ack => ct_core_CP_34_elements(154)); -- 
    -- CP-element group 155:  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	152 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_Update/cr
      -- CP-element group 155: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_update_start_
      -- CP-element group 155: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_sample_completed_
      -- 
    ra_1196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_589_inst_ack_0, ack => ct_core_CP_34_elements(155)); -- 
    cr_1200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(155), ack => RPIPE_ConvTranspose_input_pipe_589_inst_req_1); -- 
    -- CP-element group 156:  transition  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (6) 
      -- CP-element group 156: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_589_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_Sample/$entry
      -- 
    ca_1201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_589_inst_ack_1, ack => ct_core_CP_34_elements(156)); -- 
    rr_1209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(156), ack => type_cast_593_inst_req_0); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_sample_completed_
      -- 
    ra_1210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_0, ack => ct_core_CP_34_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	501 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_update_completed_
      -- 
    ca_1215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_1, ack => ct_core_CP_34_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	126 
    -- CP-element group 159: 	130 
    -- CP-element group 159: 	134 
    -- CP-element group 159: 	138 
    -- CP-element group 159: 	142 
    -- CP-element group 159: 	146 
    -- CP-element group 159: 	150 
    -- CP-element group 159: 	154 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (9) 
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/word_access_start/word_0/rr
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/word_access_start/word_0/$entry
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/word_access_start/$entry
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/ptr_deref_601_Split/split_ack
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/ptr_deref_601_Split/split_req
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/ptr_deref_601_Split/$exit
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/ptr_deref_601_Split/$entry
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_sample_start_
      -- 
    rr_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(159), ack => ptr_deref_601_store_0_req_0); -- 
    ct_core_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(126) & ct_core_CP_34_elements(130) & ct_core_CP_34_elements(134) & ct_core_CP_34_elements(138) & ct_core_CP_34_elements(142) & ct_core_CP_34_elements(146) & ct_core_CP_34_elements(150) & ct_core_CP_34_elements(154) & ct_core_CP_34_elements(158);
      gj_ct_core_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (5) 
      -- CP-element group 160: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/word_access_start/word_0/ra
      -- CP-element group 160: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/word_access_start/word_0/$exit
      -- CP-element group 160: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/word_access_start/$exit
      -- CP-element group 160: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_sample_completed_
      -- 
    ra_1254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_601_store_0_ack_0, ack => ct_core_CP_34_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	501 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (5) 
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Update/word_access_complete/word_0/ca
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Update/word_access_complete/word_0/$exit
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Update/word_access_complete/$exit
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_update_completed_
      -- 
    ca_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_601_store_0_ack_1, ack => ct_core_CP_34_elements(161)); -- 
    -- CP-element group 162:  branch  join  transition  place  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	123 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (10) 
      -- CP-element group 162: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614__exit__
      -- CP-element group 162: 	 branch_block_stmt_25/if_stmt_615__entry__
      -- CP-element group 162: 	 branch_block_stmt_25/if_stmt_615_else_link/$entry
      -- CP-element group 162: 	 branch_block_stmt_25/if_stmt_615_if_link/$entry
      -- CP-element group 162: 	 branch_block_stmt_25/if_stmt_615_dead_link/$entry
      -- CP-element group 162: 	 branch_block_stmt_25/R_exitcond2_616_place
      -- CP-element group 162: 	 branch_block_stmt_25/if_stmt_615_eval_test/branch_req
      -- CP-element group 162: 	 branch_block_stmt_25/if_stmt_615_eval_test/$exit
      -- CP-element group 162: 	 branch_block_stmt_25/if_stmt_615_eval_test/$entry
      -- CP-element group 162: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/$exit
      -- 
    branch_req_1273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(162), ack => if_stmt_615_branch_req_0); -- 
    ct_core_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(123) & ct_core_CP_34_elements(161);
      gj_ct_core_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  merge  transition  place  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	495 
    -- CP-element group 163:  members (13) 
      -- CP-element group 163: 	 branch_block_stmt_25/merge_stmt_399__exit__
      -- CP-element group 163: 	 branch_block_stmt_25/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader
      -- CP-element group 163: 	 branch_block_stmt_25/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit
      -- CP-element group 163: 	 branch_block_stmt_25/if_stmt_615_if_link/if_choice_transition
      -- CP-element group 163: 	 branch_block_stmt_25/if_stmt_615_if_link/$exit
      -- CP-element group 163: 	 branch_block_stmt_25/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader_PhiReq/$exit
      -- CP-element group 163: 	 branch_block_stmt_25/forx_xcond171x_xpreheaderx_xloopexit_forx_xcond171x_xpreheader_PhiReq/$entry
      -- CP-element group 163: 	 branch_block_stmt_25/merge_stmt_399_PhiAck/dummy
      -- CP-element group 163: 	 branch_block_stmt_25/merge_stmt_399_PhiAck/$exit
      -- CP-element group 163: 	 branch_block_stmt_25/merge_stmt_399_PhiAck/$entry
      -- CP-element group 163: 	 branch_block_stmt_25/merge_stmt_399_PhiReqMerge
      -- CP-element group 163: 	 branch_block_stmt_25/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 163: 	 branch_block_stmt_25/forx_xbody_forx_xcond171x_xpreheaderx_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_615_branch_ack_1, ack => ct_core_CP_34_elements(163)); -- 
    -- CP-element group 164:  fork  transition  place  input  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	497 
    -- CP-element group 164: 	498 
    -- CP-element group 164:  members (12) 
      -- CP-element group 164: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/SplitProtocol/Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/if_stmt_615_else_link/$exit
      -- CP-element group 164: 	 branch_block_stmt_25/forx_xbody_forx_xbody
      -- CP-element group 164: 	 branch_block_stmt_25/if_stmt_615_else_link/else_choice_transition
      -- CP-element group 164: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/SplitProtocol/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/SplitProtocol/Sample/rr
      -- CP-element group 164: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/$entry
      -- CP-element group 164: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/SplitProtocol/Update/cr
      -- CP-element group 164: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/SplitProtocol/Update/$entry
      -- 
    else_choice_transition_1282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_615_branch_ack_0, ack => ct_core_CP_34_elements(164)); -- 
    rr_3114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(164), ack => type_cast_458_inst_req_0); -- 
    cr_3119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(164), ack => type_cast_458_inst_req_1); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	119 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_Sample/ra
      -- 
    ra_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_642_inst_ack_0, ack => ct_core_CP_34_elements(165)); -- 
    -- CP-element group 166:  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	119 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	502 
    -- CP-element group 166:  members (9) 
      -- CP-element group 166: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656__exit__
      -- CP-element group 166: 	 branch_block_stmt_25/bbx_xnph465_forx_xbody177
      -- CP-element group 166: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/$exit
      -- CP-element group 166: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_Update/ca
      -- CP-element group 166: 	 branch_block_stmt_25/assign_stmt_627_to_assign_stmt_656/type_cast_642_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_25/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_25/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_659/$entry
      -- CP-element group 166: 	 branch_block_stmt_25/bbx_xnph465_forx_xbody177_PhiReq/$entry
      -- 
    ca_1301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_642_inst_ack_1, ack => ct_core_CP_34_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	507 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	206 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_final_index_sum_regn_Sample/ack
      -- CP-element group 167: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_final_index_sum_regn_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_final_index_sum_regn_sample_complete
      -- 
    ack_1330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_671_index_offset_ack_0, ack => ct_core_CP_34_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	507 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (11) 
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_final_index_sum_regn_Update/ack
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_final_index_sum_regn_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_request/req
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_request/$entry
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_offset_calculated
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_root_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_base_plus_offset/sum_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_base_plus_offset/sum_rename_req
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_base_plus_offset/$exit
      -- CP-element group 168: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_base_plus_offset/$entry
      -- 
    ack_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_671_index_offset_ack_1, ack => ct_core_CP_34_elements(168)); -- 
    req_1344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(168), ack => addr_of_672_final_reg_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_request/ack
      -- CP-element group 169: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_request/$exit
      -- CP-element group 169: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_sample_completed_
      -- 
    ack_1345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_672_final_reg_ack_0, ack => ct_core_CP_34_elements(169)); -- 
    -- CP-element group 170:  fork  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	507 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	203 
    -- CP-element group 170:  members (19) 
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_complete/ack
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_complete/$exit
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_base_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_word_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_base_address_resized
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_base_addr_resize/$entry
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_base_addr_resize/$exit
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_base_addr_resize/base_resize_req
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_base_addr_resize/base_resize_ack
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_word_addrgen/$entry
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_word_addrgen/$exit
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_word_addrgen/root_register_req
      -- CP-element group 170: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_word_addrgen/root_register_ack
      -- 
    ack_1350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_672_final_reg_ack_1, ack => ct_core_CP_34_elements(170)); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	507 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (6) 
      -- CP-element group 171: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_Update/cr
      -- CP-element group 171: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_Sample/ra
      -- CP-element group 171: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_update_start_
      -- CP-element group 171: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_sample_completed_
      -- 
    ra_1359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_675_inst_ack_0, ack => ct_core_CP_34_elements(171)); -- 
    cr_1363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(171), ack => RPIPE_ConvTranspose_input_pipe_675_inst_req_1); -- 
    -- CP-element group 172:  fork  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172: 	175 
    -- CP-element group 172:  members (9) 
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_Update/ca
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_update_completed_
      -- 
    ca_1364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_675_inst_ack_1, ack => ct_core_CP_34_elements(172)); -- 
    rr_1372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(172), ack => type_cast_679_inst_req_0); -- 
    rr_1386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(172), ack => RPIPE_ConvTranspose_input_pipe_688_inst_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_Sample/$exit
      -- 
    ra_1373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_0, ack => ct_core_CP_34_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	507 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	203 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_update_completed_
      -- 
    ca_1378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_1, ack => ct_core_CP_34_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	172 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_update_start_
      -- CP-element group 175: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_Update/cr
      -- 
    ra_1387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_688_inst_ack_0, ack => ct_core_CP_34_elements(175)); -- 
    cr_1391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(175), ack => RPIPE_ConvTranspose_input_pipe_688_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_688_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_Sample/$entry
      -- 
    ca_1392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_688_inst_ack_1, ack => ct_core_CP_34_elements(176)); -- 
    rr_1400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(176), ack => type_cast_692_inst_req_0); -- 
    rr_1414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(176), ack => RPIPE_ConvTranspose_input_pipe_706_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_sample_completed_
      -- 
    ra_1401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_692_inst_ack_0, ack => ct_core_CP_34_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	507 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	203 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_update_completed_
      -- 
    ca_1406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_692_inst_ack_1, ack => ct_core_CP_34_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_Update/cr
      -- CP-element group 179: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_update_start_
      -- CP-element group 179: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_sample_completed_
      -- 
    ra_1415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_706_inst_ack_0, ack => ct_core_CP_34_elements(179)); -- 
    cr_1419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(179), ack => RPIPE_ConvTranspose_input_pipe_706_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_706_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_Sample/rr
      -- 
    ca_1420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_706_inst_ack_1, ack => ct_core_CP_34_elements(180)); -- 
    rr_1428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(180), ack => type_cast_710_inst_req_0); -- 
    rr_1442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(180), ack => RPIPE_ConvTranspose_input_pipe_724_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_Sample/ra
      -- 
    ra_1429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_710_inst_ack_0, ack => ct_core_CP_34_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	507 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	203 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_Update/ca
      -- 
    ca_1434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_710_inst_ack_1, ack => ct_core_CP_34_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_update_start_
      -- CP-element group 183: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_Update/cr
      -- 
    ra_1443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_724_inst_ack_0, ack => ct_core_CP_34_elements(183)); -- 
    cr_1447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(183), ack => RPIPE_ConvTranspose_input_pipe_724_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_724_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_Sample/rr
      -- 
    ca_1448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_724_inst_ack_1, ack => ct_core_CP_34_elements(184)); -- 
    rr_1456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(184), ack => type_cast_728_inst_req_0); -- 
    rr_1470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(184), ack => RPIPE_ConvTranspose_input_pipe_742_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_Sample/ra
      -- 
    ra_1457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_728_inst_ack_0, ack => ct_core_CP_34_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	507 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	203 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_Update/ca
      -- 
    ca_1462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_728_inst_ack_1, ack => ct_core_CP_34_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_update_start_
      -- CP-element group 187: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_Update/cr
      -- 
    ra_1471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_742_inst_ack_0, ack => ct_core_CP_34_elements(187)); -- 
    cr_1475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(187), ack => RPIPE_ConvTranspose_input_pipe_742_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_742_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_Sample/rr
      -- 
    ca_1476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_742_inst_ack_1, ack => ct_core_CP_34_elements(188)); -- 
    rr_1484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(188), ack => type_cast_746_inst_req_0); -- 
    rr_1498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(188), ack => RPIPE_ConvTranspose_input_pipe_760_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_Sample/ra
      -- 
    ra_1485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_746_inst_ack_0, ack => ct_core_CP_34_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	507 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	203 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_Update/ca
      -- 
    ca_1490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_746_inst_ack_1, ack => ct_core_CP_34_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_update_start_
      -- CP-element group 191: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_Update/cr
      -- 
    ra_1499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_760_inst_ack_0, ack => ct_core_CP_34_elements(191)); -- 
    cr_1503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(191), ack => RPIPE_ConvTranspose_input_pipe_760_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_760_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_Sample/rr
      -- 
    ca_1504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_760_inst_ack_1, ack => ct_core_CP_34_elements(192)); -- 
    rr_1512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(192), ack => type_cast_764_inst_req_0); -- 
    rr_1526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(192), ack => RPIPE_ConvTranspose_input_pipe_778_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_Sample/ra
      -- 
    ra_1513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_0, ack => ct_core_CP_34_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	507 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	203 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_Update/ca
      -- 
    ca_1518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_1, ack => ct_core_CP_34_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_update_start_
      -- CP-element group 195: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_Update/cr
      -- 
    ra_1527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_778_inst_ack_0, ack => ct_core_CP_34_elements(195)); -- 
    cr_1531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(195), ack => RPIPE_ConvTranspose_input_pipe_778_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_778_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_Sample/rr
      -- 
    ca_1532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_778_inst_ack_1, ack => ct_core_CP_34_elements(196)); -- 
    rr_1540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(196), ack => type_cast_782_inst_req_0); -- 
    rr_1554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(196), ack => RPIPE_ConvTranspose_input_pipe_796_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_Sample/ra
      -- 
    ra_1541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_782_inst_ack_0, ack => ct_core_CP_34_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	507 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	203 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_Update/ca
      -- 
    ca_1546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_782_inst_ack_1, ack => ct_core_CP_34_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_update_start_
      -- CP-element group 199: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_Update/cr
      -- 
    ra_1555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_796_inst_ack_0, ack => ct_core_CP_34_elements(199)); -- 
    cr_1559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(199), ack => RPIPE_ConvTranspose_input_pipe_796_inst_req_1); -- 
    -- CP-element group 200:  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (6) 
      -- CP-element group 200: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_796_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_Sample/rr
      -- 
    ca_1560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_796_inst_ack_1, ack => ct_core_CP_34_elements(200)); -- 
    rr_1568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(200), ack => type_cast_800_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_Sample/ra
      -- 
    ra_1569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_800_inst_ack_0, ack => ct_core_CP_34_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	507 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_Update/ca
      -- 
    ca_1574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_800_inst_ack_1, ack => ct_core_CP_34_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	170 
    -- CP-element group 203: 	174 
    -- CP-element group 203: 	178 
    -- CP-element group 203: 	182 
    -- CP-element group 203: 	186 
    -- CP-element group 203: 	190 
    -- CP-element group 203: 	194 
    -- CP-element group 203: 	198 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (9) 
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/ptr_deref_808_Split/$entry
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/ptr_deref_808_Split/$exit
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/ptr_deref_808_Split/split_req
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/ptr_deref_808_Split/split_ack
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/word_access_start/$entry
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/word_access_start/word_0/$entry
      -- CP-element group 203: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/word_access_start/word_0/rr
      -- 
    rr_1612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(203), ack => ptr_deref_808_store_0_req_0); -- 
    ct_core_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(170) & ct_core_CP_34_elements(174) & ct_core_CP_34_elements(178) & ct_core_CP_34_elements(182) & ct_core_CP_34_elements(186) & ct_core_CP_34_elements(190) & ct_core_CP_34_elements(194) & ct_core_CP_34_elements(198) & ct_core_CP_34_elements(202);
      gj_ct_core_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (5) 
      -- CP-element group 204: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/word_access_start/$exit
      -- CP-element group 204: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/word_access_start/word_0/$exit
      -- CP-element group 204: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Sample/word_access_start/word_0/ra
      -- 
    ra_1613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_808_store_0_ack_0, ack => ct_core_CP_34_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	507 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (5) 
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Update/word_access_complete/$exit
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Update/word_access_complete/word_0/$exit
      -- CP-element group 205: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Update/word_access_complete/word_0/ca
      -- 
    ca_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_808_store_0_ack_1, ack => ct_core_CP_34_elements(205)); -- 
    -- CP-element group 206:  branch  join  transition  place  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	167 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (10) 
      -- CP-element group 206: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821__exit__
      -- CP-element group 206: 	 branch_block_stmt_25/if_stmt_822__entry__
      -- CP-element group 206: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/$exit
      -- CP-element group 206: 	 branch_block_stmt_25/if_stmt_822_dead_link/$entry
      -- CP-element group 206: 	 branch_block_stmt_25/if_stmt_822_eval_test/$entry
      -- CP-element group 206: 	 branch_block_stmt_25/if_stmt_822_eval_test/$exit
      -- CP-element group 206: 	 branch_block_stmt_25/if_stmt_822_eval_test/branch_req
      -- CP-element group 206: 	 branch_block_stmt_25/R_exitcond22_823_place
      -- CP-element group 206: 	 branch_block_stmt_25/if_stmt_822_if_link/$entry
      -- CP-element group 206: 	 branch_block_stmt_25/if_stmt_822_else_link/$entry
      -- 
    branch_req_1632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(206), ack => if_stmt_822_branch_req_0); -- 
    ct_core_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(167) & ct_core_CP_34_elements(205);
      gj_ct_core_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  merge  transition  place  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	508 
    -- CP-element group 207:  members (13) 
      -- CP-element group 207: 	 branch_block_stmt_25/merge_stmt_828__exit__
      -- CP-element group 207: 	 branch_block_stmt_25/forx_xend231x_xloopexit_forx_xend231
      -- CP-element group 207: 	 branch_block_stmt_25/merge_stmt_828_PhiAck/$exit
      -- CP-element group 207: 	 branch_block_stmt_25/merge_stmt_828_PhiAck/dummy
      -- CP-element group 207: 	 branch_block_stmt_25/forx_xend231x_xloopexit_forx_xend231_PhiReq/$exit
      -- CP-element group 207: 	 branch_block_stmt_25/forx_xbody177_forx_xend231x_xloopexit_PhiReq/$exit
      -- CP-element group 207: 	 branch_block_stmt_25/if_stmt_822_if_link/$exit
      -- CP-element group 207: 	 branch_block_stmt_25/if_stmt_822_if_link/if_choice_transition
      -- CP-element group 207: 	 branch_block_stmt_25/forx_xbody177_forx_xend231x_xloopexit
      -- CP-element group 207: 	 branch_block_stmt_25/merge_stmt_828_PhiAck/$entry
      -- CP-element group 207: 	 branch_block_stmt_25/forx_xend231x_xloopexit_forx_xend231_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_25/merge_stmt_828_PhiReqMerge
      -- CP-element group 207: 	 branch_block_stmt_25/forx_xbody177_forx_xend231x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_822_branch_ack_1, ack => ct_core_CP_34_elements(207)); -- 
    -- CP-element group 208:  fork  transition  place  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	503 
    -- CP-element group 208: 	504 
    -- CP-element group 208:  members (12) 
      -- CP-element group 208: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/SplitProtocol/Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/SplitProtocol/Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/$entry
      -- CP-element group 208: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/$entry
      -- CP-element group 208: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/SplitProtocol/$entry
      -- CP-element group 208: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/SplitProtocol/Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_25/if_stmt_822_else_link/$exit
      -- CP-element group 208: 	 branch_block_stmt_25/if_stmt_822_else_link/else_choice_transition
      -- CP-element group 208: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177
      -- CP-element group 208: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/SplitProtocol/Update/cr
      -- CP-element group 208: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/$entry
      -- CP-element group 208: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/$entry
      -- 
    else_choice_transition_1641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_822_branch_ack_0, ack => ct_core_CP_34_elements(208)); -- 
    rr_3168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(208), ack => type_cast_665_inst_req_0); -- 
    cr_3173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(208), ack => type_cast_665_inst_req_1); -- 
    -- CP-element group 209:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	508 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	211 
    -- CP-element group 209: 	212 
    -- CP-element group 209:  members (18) 
      -- CP-element group 209: 	 branch_block_stmt_25/merge_stmt_843_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_25/merge_stmt_843__exit__
      -- CP-element group 209: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878__entry__
      -- CP-element group 209: 	 branch_block_stmt_25/if_stmt_837_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_25/if_stmt_837_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_25/forx_xend250_bbx_xnph450
      -- CP-element group 209: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/$entry
      -- CP-element group 209: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_sample_start_
      -- CP-element group 209: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_update_start_
      -- CP-element group 209: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_Sample/$entry
      -- CP-element group 209: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_Sample/rr
      -- CP-element group 209: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_Update/$entry
      -- CP-element group 209: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_Update/cr
      -- CP-element group 209: 	 branch_block_stmt_25/merge_stmt_843_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_25/merge_stmt_843_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_25/merge_stmt_843_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_25/forx_xend250_bbx_xnph450_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_25/forx_xend250_bbx_xnph450_PhiReq/$entry
      -- 
    if_choice_transition_1659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_837_branch_ack_1, ack => ct_core_CP_34_elements(209)); -- 
    rr_1676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(209), ack => type_cast_864_inst_req_0); -- 
    cr_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(209), ack => type_cast_864_inst_req_1); -- 
    -- CP-element group 210:  transition  place  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	508 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	515 
    -- CP-element group 210:  members (5) 
      -- CP-element group 210: 	 branch_block_stmt_25/if_stmt_837_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_25/if_stmt_837_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xend250_forx_xend273
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_25/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_837_branch_ack_0, ack => ct_core_CP_34_elements(210)); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_Sample/ra
      -- 
    ra_1677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_864_inst_ack_0, ack => ct_core_CP_34_elements(211)); -- 
    -- CP-element group 212:  transition  place  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	209 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	509 
    -- CP-element group 212:  members (9) 
      -- CP-element group 212: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878__exit__
      -- CP-element group 212: 	 branch_block_stmt_25/bbx_xnph451_forx_xbody266
      -- CP-element group 212: 	 branch_block_stmt_25/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/$exit
      -- CP-element group 212: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_25/assign_stmt_849_to_assign_stmt_878/type_cast_864_Update/ca
      -- CP-element group 212: 	 branch_block_stmt_25/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_881/$entry
      -- CP-element group 212: 	 branch_block_stmt_25/bbx_xnph451_forx_xbody266_PhiReq/$entry
      -- 
    ca_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_864_inst_ack_1, ack => ct_core_CP_34_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	514 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	219 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_final_index_sum_regn_sample_complete
      -- CP-element group 213: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_final_index_sum_regn_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_final_index_sum_regn_Sample/ack
      -- 
    ack_1711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_893_index_offset_ack_0, ack => ct_core_CP_34_elements(213)); -- 
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	514 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (11) 
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_root_address_calculated
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_offset_calculated
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_final_index_sum_regn_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_final_index_sum_regn_Update/ack
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_base_plus_offset/$entry
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_base_plus_offset/$exit
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_base_plus_offset/sum_rename_req
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_base_plus_offset/sum_rename_ack
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_request/$entry
      -- CP-element group 214: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_request/req
      -- 
    ack_1716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_893_index_offset_ack_1, ack => ct_core_CP_34_elements(214)); -- 
    req_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(214), ack => addr_of_894_final_reg_req_0); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_request/$exit
      -- CP-element group 215: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_request/ack
      -- 
    ack_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_894_final_reg_ack_0, ack => ct_core_CP_34_elements(215)); -- 
    -- CP-element group 216:  join  fork  transition  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	514 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (28) 
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_complete/$exit
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_complete/ack
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_base_address_calculated
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_word_address_calculated
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_root_address_calculated
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_base_address_resized
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_base_addr_resize/$entry
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_base_addr_resize/$exit
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_base_addr_resize/base_resize_req
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_base_addr_resize/base_resize_ack
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_base_plus_offset/$entry
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_base_plus_offset/$exit
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_base_plus_offset/sum_rename_req
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_base_plus_offset/sum_rename_ack
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_word_addrgen/$entry
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_word_addrgen/$exit
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_word_addrgen/root_register_req
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_word_addrgen/root_register_ack
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/ptr_deref_897_Split/$entry
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/ptr_deref_897_Split/$exit
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/ptr_deref_897_Split/split_req
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/ptr_deref_897_Split/split_ack
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/word_access_start/$entry
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/word_access_start/word_0/$entry
      -- CP-element group 216: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/word_access_start/word_0/rr
      -- 
    ack_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_894_final_reg_ack_1, ack => ct_core_CP_34_elements(216)); -- 
    rr_1769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(216), ack => ptr_deref_897_store_0_req_0); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (5) 
      -- CP-element group 217: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/word_access_start/$exit
      -- CP-element group 217: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/word_access_start/word_0/$exit
      -- CP-element group 217: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Sample/word_access_start/word_0/ra
      -- 
    ra_1770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_897_store_0_ack_0, ack => ct_core_CP_34_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	514 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (5) 
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Update/word_access_complete/$exit
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Update/word_access_complete/word_0/$exit
      -- CP-element group 218: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Update/word_access_complete/word_0/ca
      -- 
    ca_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_897_store_0_ack_1, ack => ct_core_CP_34_elements(218)); -- 
    -- CP-element group 219:  branch  join  transition  place  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: 	213 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (10) 
      -- CP-element group 219: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911__exit__
      -- CP-element group 219: 	 branch_block_stmt_25/if_stmt_912__entry__
      -- CP-element group 219: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/$exit
      -- CP-element group 219: 	 branch_block_stmt_25/if_stmt_912_dead_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_25/if_stmt_912_eval_test/$entry
      -- CP-element group 219: 	 branch_block_stmt_25/if_stmt_912_eval_test/$exit
      -- CP-element group 219: 	 branch_block_stmt_25/if_stmt_912_eval_test/branch_req
      -- CP-element group 219: 	 branch_block_stmt_25/R_exitcond_913_place
      -- CP-element group 219: 	 branch_block_stmt_25/if_stmt_912_if_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_25/if_stmt_912_else_link/$entry
      -- 
    branch_req_1789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(219), ack => if_stmt_912_branch_req_0); -- 
    ct_core_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(218) & ct_core_CP_34_elements(213);
      gj_ct_core_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  merge  transition  place  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	515 
    -- CP-element group 220:  members (13) 
      -- CP-element group 220: 	 branch_block_stmt_25/merge_stmt_918__exit__
      -- CP-element group 220: 	 branch_block_stmt_25/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 220: 	 branch_block_stmt_25/if_stmt_912_if_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_25/if_stmt_912_if_link/if_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_25/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 220: 	 branch_block_stmt_25/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_25/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 220: 	 branch_block_stmt_25/merge_stmt_918_PhiReqMerge
      -- CP-element group 220: 	 branch_block_stmt_25/merge_stmt_918_PhiAck/$entry
      -- CP-element group 220: 	 branch_block_stmt_25/merge_stmt_918_PhiAck/$exit
      -- CP-element group 220: 	 branch_block_stmt_25/merge_stmt_918_PhiAck/dummy
      -- CP-element group 220: 	 branch_block_stmt_25/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_25/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_912_branch_ack_1, ack => ct_core_CP_34_elements(220)); -- 
    -- CP-element group 221:  fork  transition  place  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	510 
    -- CP-element group 221: 	511 
    -- CP-element group 221:  members (12) 
      -- CP-element group 221: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/$entry
      -- CP-element group 221: 	 branch_block_stmt_25/if_stmt_912_else_link/$exit
      -- CP-element group 221: 	 branch_block_stmt_25/if_stmt_912_else_link/else_choice_transition
      -- CP-element group 221: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/SplitProtocol/Update/cr
      -- CP-element group 221: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/$entry
      -- CP-element group 221: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/SplitProtocol/Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/SplitProtocol/Sample/rr
      -- CP-element group 221: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/SplitProtocol/Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/SplitProtocol/$entry
      -- CP-element group 221: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/$entry
      -- 
    else_choice_transition_1798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_912_branch_ack_0, ack => ct_core_CP_34_elements(221)); -- 
    cr_3250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(221), ack => type_cast_887_inst_req_1); -- 
    rr_3245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(221), ack => type_cast_887_inst_req_0); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	515 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_sample_completed_
      -- CP-element group 222: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_Sample/cra
      -- 
    cra_1812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_923_call_ack_0, ack => ct_core_CP_34_elements(222)); -- 
    -- CP-element group 223:  transition  place  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	515 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (10) 
      -- CP-element group 223: 	 branch_block_stmt_25/call_stmt_923__exit__
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_928_to_assign_stmt_955__entry__
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_928_to_assign_stmt_955__exit__
      -- CP-element group 223: 	 branch_block_stmt_25/do_while_stmt_956__entry__
      -- CP-element group 223: 	 branch_block_stmt_25/call_stmt_923/$exit
      -- CP-element group 223: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_update_completed_
      -- CP-element group 223: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_Update/cca
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_928_to_assign_stmt_955/$entry
      -- CP-element group 223: 	 branch_block_stmt_25/assign_stmt_928_to_assign_stmt_955/$exit
      -- 
    cca_1817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_923_call_ack_1, ack => ct_core_CP_34_elements(223)); -- 
    -- CP-element group 224:  transition  place  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	230 
    -- CP-element group 224:  members (2) 
      -- CP-element group 224: 	 branch_block_stmt_25/do_while_stmt_956/$entry
      -- CP-element group 224: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956__entry__
      -- 
    ct_core_CP_34_elements(224) <= ct_core_CP_34_elements(223);
    -- CP-element group 225:  merge  place  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	396 
    -- CP-element group 225:  members (1) 
      -- CP-element group 225: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956__exit__
      -- 
    -- Element group ct_core_CP_34_elements(225) is bound as output of CP function.
    -- CP-element group 226:  merge  place  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	229 
    -- CP-element group 226:  members (1) 
      -- CP-element group 226: 	 branch_block_stmt_25/do_while_stmt_956/loop_back
      -- 
    -- Element group ct_core_CP_34_elements(226) is bound as output of CP function.
    -- CP-element group 227:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	232 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	394 
    -- CP-element group 227: 	395 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_25/do_while_stmt_956/condition_done
      -- CP-element group 227: 	 branch_block_stmt_25/do_while_stmt_956/loop_exit/$entry
      -- CP-element group 227: 	 branch_block_stmt_25/do_while_stmt_956/loop_taken/$entry
      -- 
    ct_core_CP_34_elements(227) <= ct_core_CP_34_elements(232);
    -- CP-element group 228:  branch  place  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	393 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (1) 
      -- CP-element group 228: 	 branch_block_stmt_25/do_while_stmt_956/loop_body_done
      -- 
    ct_core_CP_34_elements(228) <= ct_core_CP_34_elements(393);
    -- CP-element group 229:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	226 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	241 
    -- CP-element group 229: 	260 
    -- CP-element group 229: 	279 
    -- CP-element group 229: 	298 
    -- CP-element group 229: 	317 
    -- CP-element group 229: 	336 
    -- CP-element group 229:  members (1) 
      -- CP-element group 229: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/back_edge_to_loop_body
      -- 
    ct_core_CP_34_elements(229) <= ct_core_CP_34_elements(226);
    -- CP-element group 230:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	224 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	243 
    -- CP-element group 230: 	262 
    -- CP-element group 230: 	281 
    -- CP-element group 230: 	300 
    -- CP-element group 230: 	319 
    -- CP-element group 230: 	338 
    -- CP-element group 230:  members (1) 
      -- CP-element group 230: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/first_time_through_loop_body
      -- 
    ct_core_CP_34_elements(230) <= ct_core_CP_34_elements(224);
    -- CP-element group 231:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	237 
    -- CP-element group 231: 	238 
    -- CP-element group 231: 	254 
    -- CP-element group 231: 	255 
    -- CP-element group 231: 	273 
    -- CP-element group 231: 	274 
    -- CP-element group 231: 	292 
    -- CP-element group 231: 	293 
    -- CP-element group 231: 	311 
    -- CP-element group 231: 	312 
    -- CP-element group 231: 	361 
    -- CP-element group 231: 	363 
    -- CP-element group 231: 	376 
    -- CP-element group 231: 	380 
    -- CP-element group 231: 	384 
    -- CP-element group 231: 	388 
    -- CP-element group 231: 	392 
    -- CP-element group 231: 	330 
    -- CP-element group 231: 	331 
    -- CP-element group 231: 	350 
    -- CP-element group 231: 	351 
    -- CP-element group 231:  members (2) 
      -- CP-element group 231: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/$entry
      -- CP-element group 231: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/loop_body_start
      -- 
    -- Element group ct_core_CP_34_elements(231) is bound as output of CP function.
    -- CP-element group 232:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	236 
    -- CP-element group 232: 	240 
    -- CP-element group 232: 	259 
    -- CP-element group 232: 	278 
    -- CP-element group 232: 	379 
    -- CP-element group 232: 	383 
    -- CP-element group 232: 	391 
    -- CP-element group 232: 	392 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	227 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/condition_evaluated
      -- 
    condition_evaluated_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(232), ack => do_while_stmt_956_branch_req_0); -- 
    ct_core_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(236) & ct_core_CP_34_elements(240) & ct_core_CP_34_elements(259) & ct_core_CP_34_elements(278) & ct_core_CP_34_elements(379) & ct_core_CP_34_elements(383) & ct_core_CP_34_elements(391) & ct_core_CP_34_elements(392);
      gj_ct_core_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	237 
    -- CP-element group 233: 	254 
    -- CP-element group 233: 	273 
    -- CP-element group 233: 	292 
    -- CP-element group 233: 	311 
    -- CP-element group 233: 	330 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	236 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	256 
    -- CP-element group 233: 	275 
    -- CP-element group 233: 	294 
    -- CP-element group 233: 	313 
    -- CP-element group 233: 	332 
    -- CP-element group 233:  members (2) 
      -- CP-element group 233: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/aggregated_phi_sample_req
      -- CP-element group 233: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_sample_start__ps
      -- 
    ct_core_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(237) & ct_core_CP_34_elements(254) & ct_core_CP_34_elements(273) & ct_core_CP_34_elements(292) & ct_core_CP_34_elements(311) & ct_core_CP_34_elements(330) & ct_core_CP_34_elements(236);
      gj_ct_core_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	239 
    -- CP-element group 234: 	257 
    -- CP-element group 234: 	276 
    -- CP-element group 234: 	295 
    -- CP-element group 234: 	314 
    -- CP-element group 234: 	333 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	377 
    -- CP-element group 234: 	381 
    -- CP-element group 234: 	385 
    -- CP-element group 234: 	393 
    -- CP-element group 234: marked-successors 
    -- CP-element group 234: 	237 
    -- CP-element group 234: 	254 
    -- CP-element group 234: 	273 
    -- CP-element group 234: 	292 
    -- CP-element group 234: 	311 
    -- CP-element group 234: 	330 
    -- CP-element group 234:  members (7) 
      -- CP-element group 234: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/aggregated_phi_sample_ack
      -- CP-element group 234: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_sample_completed_
      -- 
    ct_core_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(239) & ct_core_CP_34_elements(257) & ct_core_CP_34_elements(276) & ct_core_CP_34_elements(295) & ct_core_CP_34_elements(314) & ct_core_CP_34_elements(333);
      gj_ct_core_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	238 
    -- CP-element group 235: 	255 
    -- CP-element group 235: 	274 
    -- CP-element group 235: 	293 
    -- CP-element group 235: 	312 
    -- CP-element group 235: 	331 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	258 
    -- CP-element group 235: 	277 
    -- CP-element group 235: 	296 
    -- CP-element group 235: 	315 
    -- CP-element group 235: 	334 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/aggregated_phi_update_req
      -- CP-element group 235: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_update_start__ps
      -- 
    ct_core_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(238) & ct_core_CP_34_elements(255) & ct_core_CP_34_elements(274) & ct_core_CP_34_elements(293) & ct_core_CP_34_elements(312) & ct_core_CP_34_elements(331);
      gj_ct_core_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	240 
    -- CP-element group 236: 	259 
    -- CP-element group 236: 	278 
    -- CP-element group 236: 	297 
    -- CP-element group 236: 	316 
    -- CP-element group 236: 	335 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	232 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	233 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/aggregated_phi_update_ack
      -- 
    ct_core_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(240) & ct_core_CP_34_elements(259) & ct_core_CP_34_elements(278) & ct_core_CP_34_elements(297) & ct_core_CP_34_elements(316) & ct_core_CP_34_elements(335);
      gj_ct_core_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  join  transition  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	231 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	234 
    -- CP-element group 237: 	379 
    -- CP-element group 237: 	383 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	233 
    -- CP-element group 237:  members (1) 
      -- CP-element group 237: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_sample_start_
      -- 
    ct_core_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(234) & ct_core_CP_34_elements(379) & ct_core_CP_34_elements(383);
      gj_ct_core_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  join  transition  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	231 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	235 
    -- CP-element group 238:  members (1) 
      -- CP-element group 238: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_update_start_
      -- 
    ct_core_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(240);
      gj_ct_core_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  join  transition  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	234 
    -- CP-element group 239:  members (1) 
      -- CP-element group 239: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_sample_completed__ps
      -- 
    -- Element group ct_core_CP_34_elements(239) is bound as output of CP function.
    -- CP-element group 240:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	232 
    -- CP-element group 240: 	236 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	238 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_update_completed__ps
      -- 
    -- Element group ct_core_CP_34_elements(240) is bound as output of CP function.
    -- CP-element group 241:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	229 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (1) 
      -- CP-element group 241: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_loopback_trigger
      -- 
    ct_core_CP_34_elements(241) <= ct_core_CP_34_elements(229);
    -- CP-element group 242:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: successors 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_loopback_sample_req
      -- CP-element group 242: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_loopback_sample_req_ps
      -- 
    phi_stmt_958_loopback_sample_req_1850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_958_loopback_sample_req_1850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(242), ack => phi_stmt_958_req_1); -- 
    -- Element group ct_core_CP_34_elements(242) is bound as output of CP function.
    -- CP-element group 243:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	230 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (1) 
      -- CP-element group 243: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_entry_trigger
      -- 
    ct_core_CP_34_elements(243) <= ct_core_CP_34_elements(230);
    -- CP-element group 244:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (2) 
      -- CP-element group 244: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_entry_sample_req
      -- CP-element group 244: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_entry_sample_req_ps
      -- 
    phi_stmt_958_entry_sample_req_1853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_958_entry_sample_req_1853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(244), ack => phi_stmt_958_req_0); -- 
    -- Element group ct_core_CP_34_elements(244) is bound as output of CP function.
    -- CP-element group 245:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: successors 
    -- CP-element group 245:  members (2) 
      -- CP-element group 245: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_phi_mux_ack
      -- CP-element group 245: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_958_phi_mux_ack_ps
      -- 
    phi_stmt_958_phi_mux_ack_1856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_958_ack_0, ack => ct_core_CP_34_elements(245)); -- 
    -- CP-element group 246:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (4) 
      -- CP-element group 246: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim0_init_960_sample_start__ps
      -- CP-element group 246: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim0_init_960_sample_completed__ps
      -- CP-element group 246: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim0_init_960_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim0_init_960_sample_completed_
      -- 
    -- Element group ct_core_CP_34_elements(246) is bound as output of CP function.
    -- CP-element group 247:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	249 
    -- CP-element group 247:  members (2) 
      -- CP-element group 247: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim0_init_960_update_start__ps
      -- CP-element group 247: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim0_init_960_update_start_
      -- 
    -- Element group ct_core_CP_34_elements(247) is bound as output of CP function.
    -- CP-element group 248:  join  transition  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	249 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (1) 
      -- CP-element group 248: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim0_init_960_update_completed__ps
      -- 
    ct_core_CP_34_elements(248) <= ct_core_CP_34_elements(249);
    -- CP-element group 249:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	248 
    -- CP-element group 249:  members (1) 
      -- CP-element group 249: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim0_init_960_update_completed_
      -- 
    -- Element group ct_core_CP_34_elements(249) is a control-delay.
    cp_element_249_delay: control_delay_element  generic map(name => " 249_delay", delay_value => 1)  port map(req => ct_core_CP_34_elements(247), ack => ct_core_CP_34_elements(249), clk => clk, reset =>reset);
    -- CP-element group 250:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (4) 
      -- CP-element group 250: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_sample_start__ps
      -- CP-element group 250: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_Sample/req
      -- 
    req_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(250), ack => next_input_dim0_1149_961_buf_req_0); -- 
    -- Element group ct_core_CP_34_elements(250) is bound as output of CP function.
    -- CP-element group 251:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	253 
    -- CP-element group 251:  members (4) 
      -- CP-element group 251: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_update_start__ps
      -- CP-element group 251: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_update_start_
      -- CP-element group 251: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_Update/req
      -- 
    req_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(251), ack => next_input_dim0_1149_961_buf_req_1); -- 
    -- Element group ct_core_CP_34_elements(251) is bound as output of CP function.
    -- CP-element group 252:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252:  members (4) 
      -- CP-element group 252: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_sample_completed__ps
      -- CP-element group 252: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_Sample/ack
      -- 
    ack_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim0_1149_961_buf_ack_0, ack => ct_core_CP_34_elements(252)); -- 
    -- CP-element group 253:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	251 
    -- CP-element group 253: successors 
    -- CP-element group 253:  members (4) 
      -- CP-element group 253: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_update_completed__ps
      -- CP-element group 253: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim0_961_Update/ack
      -- 
    ack_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim0_1149_961_buf_ack_1, ack => ct_core_CP_34_elements(253)); -- 
    -- CP-element group 254:  join  transition  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	231 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	234 
    -- CP-element group 254: 	379 
    -- CP-element group 254: 	383 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	233 
    -- CP-element group 254:  members (1) 
      -- CP-element group 254: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_sample_start_
      -- 
    ct_core_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(234) & ct_core_CP_34_elements(379) & ct_core_CP_34_elements(383);
      gj_ct_core_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  join  transition  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	231 
    -- CP-element group 255: marked-predecessors 
    -- CP-element group 255: 	259 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	235 
    -- CP-element group 255:  members (1) 
      -- CP-element group 255: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_update_start_
      -- 
    ct_core_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(259);
      gj_ct_core_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	233 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (1) 
      -- CP-element group 256: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_sample_start__ps
      -- 
    ct_core_CP_34_elements(256) <= ct_core_CP_34_elements(233);
    -- CP-element group 257:  join  transition  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	234 
    -- CP-element group 257:  members (1) 
      -- CP-element group 257: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_sample_completed__ps
      -- 
    -- Element group ct_core_CP_34_elements(257) is bound as output of CP function.
    -- CP-element group 258:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	235 
    -- CP-element group 258: successors 
    -- CP-element group 258:  members (1) 
      -- CP-element group 258: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_update_start__ps
      -- 
    ct_core_CP_34_elements(258) <= ct_core_CP_34_elements(235);
    -- CP-element group 259:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	232 
    -- CP-element group 259: 	236 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	255 
    -- CP-element group 259:  members (2) 
      -- CP-element group 259: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_update_completed_
      -- CP-element group 259: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_update_completed__ps
      -- 
    -- Element group ct_core_CP_34_elements(259) is bound as output of CP function.
    -- CP-element group 260:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	229 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (1) 
      -- CP-element group 260: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_loopback_trigger
      -- 
    ct_core_CP_34_elements(260) <= ct_core_CP_34_elements(229);
    -- CP-element group 261:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: successors 
    -- CP-element group 261:  members (2) 
      -- CP-element group 261: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_loopback_sample_req
      -- CP-element group 261: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_loopback_sample_req_ps
      -- 
    phi_stmt_962_loopback_sample_req_1894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_962_loopback_sample_req_1894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(261), ack => phi_stmt_962_req_1); -- 
    -- Element group ct_core_CP_34_elements(261) is bound as output of CP function.
    -- CP-element group 262:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	230 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (1) 
      -- CP-element group 262: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_entry_trigger
      -- 
    ct_core_CP_34_elements(262) <= ct_core_CP_34_elements(230);
    -- CP-element group 263:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (2) 
      -- CP-element group 263: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_entry_sample_req
      -- CP-element group 263: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_entry_sample_req_ps
      -- 
    phi_stmt_962_entry_sample_req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_962_entry_sample_req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(263), ack => phi_stmt_962_req_0); -- 
    -- Element group ct_core_CP_34_elements(263) is bound as output of CP function.
    -- CP-element group 264:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: successors 
    -- CP-element group 264:  members (2) 
      -- CP-element group 264: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_phi_mux_ack
      -- CP-element group 264: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_962_phi_mux_ack_ps
      -- 
    phi_stmt_962_phi_mux_ack_1900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_962_ack_0, ack => ct_core_CP_34_elements(264)); -- 
    -- CP-element group 265:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (4) 
      -- CP-element group 265: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim1_init_964_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim1_init_964_sample_start__ps
      -- CP-element group 265: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim1_init_964_sample_completed__ps
      -- CP-element group 265: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim1_init_964_sample_start_
      -- 
    -- Element group ct_core_CP_34_elements(265) is bound as output of CP function.
    -- CP-element group 266:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (2) 
      -- CP-element group 266: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim1_init_964_update_start_
      -- CP-element group 266: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim1_init_964_update_start__ps
      -- 
    -- Element group ct_core_CP_34_elements(266) is bound as output of CP function.
    -- CP-element group 267:  join  transition  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	268 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (1) 
      -- CP-element group 267: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim1_init_964_update_completed__ps
      -- 
    ct_core_CP_34_elements(267) <= ct_core_CP_34_elements(268);
    -- CP-element group 268:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	267 
    -- CP-element group 268:  members (1) 
      -- CP-element group 268: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim1_init_964_update_completed_
      -- 
    -- Element group ct_core_CP_34_elements(268) is a control-delay.
    cp_element_268_delay: control_delay_element  generic map(name => " 268_delay", delay_value => 1)  port map(req => ct_core_CP_34_elements(266), ack => ct_core_CP_34_elements(268), clk => clk, reset =>reset);
    -- CP-element group 269:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (4) 
      -- CP-element group 269: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_sample_start__ps
      -- CP-element group 269: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_Sample/req
      -- 
    req_1921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(269), ack => next_input_dim1_1143_965_buf_req_0); -- 
    -- Element group ct_core_CP_34_elements(269) is bound as output of CP function.
    -- CP-element group 270:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (4) 
      -- CP-element group 270: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_update_start__ps
      -- CP-element group 270: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_Update/req
      -- CP-element group 270: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_update_start_
      -- CP-element group 270: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_Update/$entry
      -- 
    req_1926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(270), ack => next_input_dim1_1143_965_buf_req_1); -- 
    -- Element group ct_core_CP_34_elements(270) is bound as output of CP function.
    -- CP-element group 271:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271:  members (4) 
      -- CP-element group 271: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_sample_completed__ps
      -- CP-element group 271: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_sample_completed_
      -- 
    ack_1922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim1_1143_965_buf_ack_0, ack => ct_core_CP_34_elements(271)); -- 
    -- CP-element group 272:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (4) 
      -- CP-element group 272: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_update_completed__ps
      -- CP-element group 272: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim1_965_Update/ack
      -- 
    ack_1927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim1_1143_965_buf_ack_1, ack => ct_core_CP_34_elements(272)); -- 
    -- CP-element group 273:  join  transition  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	231 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	234 
    -- CP-element group 273: 	379 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	233 
    -- CP-element group 273:  members (1) 
      -- CP-element group 273: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_sample_start_
      -- 
    ct_core_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(234) & ct_core_CP_34_elements(379);
      gj_ct_core_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  join  transition  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	231 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	278 
    -- CP-element group 274: 	364 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	235 
    -- CP-element group 274:  members (1) 
      -- CP-element group 274: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_update_start_
      -- 
    ct_core_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(278) & ct_core_CP_34_elements(364);
      gj_ct_core_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	233 
    -- CP-element group 275: successors 
    -- CP-element group 275:  members (1) 
      -- CP-element group 275: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_sample_start__ps
      -- 
    ct_core_CP_34_elements(275) <= ct_core_CP_34_elements(233);
    -- CP-element group 276:  join  transition  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	234 
    -- CP-element group 276:  members (1) 
      -- CP-element group 276: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_sample_completed__ps
      -- 
    -- Element group ct_core_CP_34_elements(276) is bound as output of CP function.
    -- CP-element group 277:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	235 
    -- CP-element group 277: successors 
    -- CP-element group 277:  members (1) 
      -- CP-element group 277: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_update_start__ps
      -- 
    ct_core_CP_34_elements(277) <= ct_core_CP_34_elements(235);
    -- CP-element group 278:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	232 
    -- CP-element group 278: 	236 
    -- CP-element group 278: 	362 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	274 
    -- CP-element group 278:  members (2) 
      -- CP-element group 278: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_update_completed__ps
      -- 
    -- Element group ct_core_CP_34_elements(278) is bound as output of CP function.
    -- CP-element group 279:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	229 
    -- CP-element group 279: successors 
    -- CP-element group 279:  members (1) 
      -- CP-element group 279: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_loopback_trigger
      -- 
    ct_core_CP_34_elements(279) <= ct_core_CP_34_elements(229);
    -- CP-element group 280:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: successors 
    -- CP-element group 280:  members (2) 
      -- CP-element group 280: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_loopback_sample_req_ps
      -- CP-element group 280: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_loopback_sample_req
      -- 
    phi_stmt_966_loopback_sample_req_1938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_966_loopback_sample_req_1938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(280), ack => phi_stmt_966_req_1); -- 
    -- Element group ct_core_CP_34_elements(280) is bound as output of CP function.
    -- CP-element group 281:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	230 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (1) 
      -- CP-element group 281: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_entry_trigger
      -- 
    ct_core_CP_34_elements(281) <= ct_core_CP_34_elements(230);
    -- CP-element group 282:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: successors 
    -- CP-element group 282:  members (2) 
      -- CP-element group 282: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_entry_sample_req_ps
      -- CP-element group 282: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_entry_sample_req
      -- 
    phi_stmt_966_entry_sample_req_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_966_entry_sample_req_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(282), ack => phi_stmt_966_req_0); -- 
    -- Element group ct_core_CP_34_elements(282) is bound as output of CP function.
    -- CP-element group 283:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (2) 
      -- CP-element group 283: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_phi_mux_ack_ps
      -- CP-element group 283: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_966_phi_mux_ack
      -- 
    phi_stmt_966_phi_mux_ack_1944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_966_ack_0, ack => ct_core_CP_34_elements(283)); -- 
    -- CP-element group 284:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: successors 
    -- CP-element group 284:  members (4) 
      -- CP-element group 284: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim2_init_968_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim2_init_968_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim2_init_968_sample_completed__ps
      -- CP-element group 284: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim2_init_968_sample_start__ps
      -- 
    -- Element group ct_core_CP_34_elements(284) is bound as output of CP function.
    -- CP-element group 285:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (2) 
      -- CP-element group 285: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim2_init_968_update_start_
      -- CP-element group 285: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim2_init_968_update_start__ps
      -- 
    -- Element group ct_core_CP_34_elements(285) is bound as output of CP function.
    -- CP-element group 286:  join  transition  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	287 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (1) 
      -- CP-element group 286: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim2_init_968_update_completed__ps
      -- 
    ct_core_CP_34_elements(286) <= ct_core_CP_34_elements(287);
    -- CP-element group 287:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	286 
    -- CP-element group 287:  members (1) 
      -- CP-element group 287: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_input_dim2_init_968_update_completed_
      -- 
    -- Element group ct_core_CP_34_elements(287) is a control-delay.
    cp_element_287_delay: control_delay_element  generic map(name => " 287_delay", delay_value => 1)  port map(req => ct_core_CP_34_elements(285), ack => ct_core_CP_34_elements(287), clk => clk, reset =>reset);
    -- CP-element group 288:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (4) 
      -- CP-element group 288: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_sample_start__ps
      -- CP-element group 288: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_Sample/req
      -- 
    req_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(288), ack => next_input_dim2_1133_969_buf_req_0); -- 
    -- Element group ct_core_CP_34_elements(288) is bound as output of CP function.
    -- CP-element group 289:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (4) 
      -- CP-element group 289: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_Update/req
      -- CP-element group 289: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_update_start_
      -- CP-element group 289: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_update_start__ps
      -- CP-element group 289: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_Update/$entry
      -- 
    req_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(289), ack => next_input_dim2_1133_969_buf_req_1); -- 
    -- Element group ct_core_CP_34_elements(289) is bound as output of CP function.
    -- CP-element group 290:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: successors 
    -- CP-element group 290:  members (4) 
      -- CP-element group 290: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_sample_completed__ps
      -- CP-element group 290: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_sample_completed_
      -- CP-element group 290: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_Sample/$exit
      -- CP-element group 290: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_Sample/ack
      -- 
    ack_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim2_1133_969_buf_ack_0, ack => ct_core_CP_34_elements(290)); -- 
    -- CP-element group 291:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291:  members (4) 
      -- CP-element group 291: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_update_completed_
      -- CP-element group 291: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_update_completed__ps
      -- CP-element group 291: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_Update/ack
      -- CP-element group 291: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_input_dim2_969_Update/$exit
      -- 
    ack_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_input_dim2_1133_969_buf_ack_1, ack => ct_core_CP_34_elements(291)); -- 
    -- CP-element group 292:  join  transition  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	231 
    -- CP-element group 292: marked-predecessors 
    -- CP-element group 292: 	234 
    -- CP-element group 292: 	379 
    -- CP-element group 292: 	383 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	233 
    -- CP-element group 292:  members (1) 
      -- CP-element group 292: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_sample_start_
      -- 
    ct_core_cp_element_group_292: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_292"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(234) & ct_core_CP_34_elements(379) & ct_core_CP_34_elements(383);
      gj_ct_core_cp_element_group_292 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(292), clk => clk, reset => reset); --
    end block;
    -- CP-element group 293:  join  transition  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	231 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	297 
    -- CP-element group 293: 	364 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	235 
    -- CP-element group 293:  members (1) 
      -- CP-element group 293: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_update_start_
      -- 
    ct_core_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(297) & ct_core_CP_34_elements(364);
      gj_ct_core_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	233 
    -- CP-element group 294: successors 
    -- CP-element group 294:  members (1) 
      -- CP-element group 294: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_sample_start__ps
      -- 
    ct_core_CP_34_elements(294) <= ct_core_CP_34_elements(233);
    -- CP-element group 295:  join  transition  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	234 
    -- CP-element group 295:  members (1) 
      -- CP-element group 295: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_sample_completed__ps
      -- 
    -- Element group ct_core_CP_34_elements(295) is bound as output of CP function.
    -- CP-element group 296:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	235 
    -- CP-element group 296: successors 
    -- CP-element group 296:  members (1) 
      -- CP-element group 296: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_update_start__ps
      -- 
    ct_core_CP_34_elements(296) <= ct_core_CP_34_elements(235);
    -- CP-element group 297:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	236 
    -- CP-element group 297: 	362 
    -- CP-element group 297: marked-successors 
    -- CP-element group 297: 	293 
    -- CP-element group 297:  members (2) 
      -- CP-element group 297: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_update_completed__ps
      -- CP-element group 297: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_update_completed_
      -- 
    -- Element group ct_core_CP_34_elements(297) is bound as output of CP function.
    -- CP-element group 298:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	229 
    -- CP-element group 298: successors 
    -- CP-element group 298:  members (1) 
      -- CP-element group 298: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_loopback_trigger
      -- 
    ct_core_CP_34_elements(298) <= ct_core_CP_34_elements(229);
    -- CP-element group 299:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: successors 
    -- CP-element group 299:  members (2) 
      -- CP-element group 299: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_loopback_sample_req_ps
      -- CP-element group 299: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_loopback_sample_req
      -- 
    phi_stmt_970_loopback_sample_req_1982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_970_loopback_sample_req_1982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(299), ack => phi_stmt_970_req_1); -- 
    -- Element group ct_core_CP_34_elements(299) is bound as output of CP function.
    -- CP-element group 300:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	230 
    -- CP-element group 300: successors 
    -- CP-element group 300:  members (1) 
      -- CP-element group 300: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_entry_trigger
      -- 
    ct_core_CP_34_elements(300) <= ct_core_CP_34_elements(230);
    -- CP-element group 301:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: successors 
    -- CP-element group 301:  members (2) 
      -- CP-element group 301: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_entry_sample_req_ps
      -- CP-element group 301: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_entry_sample_req
      -- 
    phi_stmt_970_entry_sample_req_1985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_970_entry_sample_req_1985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(301), ack => phi_stmt_970_req_0); -- 
    -- Element group ct_core_CP_34_elements(301) is bound as output of CP function.
    -- CP-element group 302:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: successors 
    -- CP-element group 302:  members (2) 
      -- CP-element group 302: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_phi_mux_ack_ps
      -- CP-element group 302: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_970_phi_mux_ack
      -- 
    phi_stmt_970_phi_mux_ack_1988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_970_ack_0, ack => ct_core_CP_34_elements(302)); -- 
    -- CP-element group 303:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	305 
    -- CP-element group 303:  members (4) 
      -- CP-element group 303: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_Sample/req
      -- CP-element group 303: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_sample_start__ps
      -- 
    req_2001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(303), ack => add_dest_dim0_init_946_972_buf_req_0); -- 
    -- Element group ct_core_CP_34_elements(303) is bound as output of CP function.
    -- CP-element group 304:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	306 
    -- CP-element group 304:  members (4) 
      -- CP-element group 304: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_Update/req
      -- CP-element group 304: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_update_start__ps
      -- CP-element group 304: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_update_start_
      -- CP-element group 304: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_Update/$entry
      -- 
    req_2006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(304), ack => add_dest_dim0_init_946_972_buf_req_1); -- 
    -- Element group ct_core_CP_34_elements(304) is bound as output of CP function.
    -- CP-element group 305:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	303 
    -- CP-element group 305: successors 
    -- CP-element group 305:  members (4) 
      -- CP-element group 305: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_sample_completed__ps
      -- CP-element group 305: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_Sample/ack
      -- 
    ack_2002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim0_init_946_972_buf_ack_0, ack => ct_core_CP_34_elements(305)); -- 
    -- CP-element group 306:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	304 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (4) 
      -- CP-element group 306: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_update_completed__ps
      -- CP-element group 306: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim0_init_972_Update/$exit
      -- 
    ack_2007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim0_init_946_972_buf_ack_1, ack => ct_core_CP_34_elements(306)); -- 
    -- CP-element group 307:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	309 
    -- CP-element group 307:  members (4) 
      -- CP-element group 307: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_sample_start__ps
      -- CP-element group 307: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_sample_start_
      -- CP-element group 307: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_Sample/req
      -- CP-element group 307: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_Sample/$entry
      -- 
    req_2019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(307), ack => next_add_dest_dim0_1127_973_buf_req_0); -- 
    -- Element group ct_core_CP_34_elements(307) is bound as output of CP function.
    -- CP-element group 308:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	310 
    -- CP-element group 308:  members (4) 
      -- CP-element group 308: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_update_start__ps
      -- CP-element group 308: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_update_start_
      -- CP-element group 308: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_Update/req
      -- CP-element group 308: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_Update/$entry
      -- 
    req_2024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(308), ack => next_add_dest_dim0_1127_973_buf_req_1); -- 
    -- Element group ct_core_CP_34_elements(308) is bound as output of CP function.
    -- CP-element group 309:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	307 
    -- CP-element group 309: successors 
    -- CP-element group 309:  members (4) 
      -- CP-element group 309: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_sample_completed__ps
      -- CP-element group 309: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_Sample/$exit
      -- 
    ack_2020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim0_1127_973_buf_ack_0, ack => ct_core_CP_34_elements(309)); -- 
    -- CP-element group 310:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	308 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (4) 
      -- CP-element group 310: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_update_completed__ps
      -- CP-element group 310: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim0_973_update_completed_
      -- 
    ack_2025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim0_1127_973_buf_ack_1, ack => ct_core_CP_34_elements(310)); -- 
    -- CP-element group 311:  join  transition  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	231 
    -- CP-element group 311: marked-predecessors 
    -- CP-element group 311: 	234 
    -- CP-element group 311: 	379 
    -- CP-element group 311: 	383 
    -- CP-element group 311: 	387 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	233 
    -- CP-element group 311:  members (1) 
      -- CP-element group 311: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_sample_start_
      -- 
    ct_core_cp_element_group_311: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_311"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(234) & ct_core_CP_34_elements(379) & ct_core_CP_34_elements(383) & ct_core_CP_34_elements(387);
      gj_ct_core_cp_element_group_311 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(311), clk => clk, reset => reset); --
    end block;
    -- CP-element group 312:  join  transition  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	231 
    -- CP-element group 312: marked-predecessors 
    -- CP-element group 312: 	316 
    -- CP-element group 312: 	364 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	235 
    -- CP-element group 312:  members (1) 
      -- CP-element group 312: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_update_start_
      -- 
    ct_core_cp_element_group_312: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_312"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(316) & ct_core_CP_34_elements(364);
      gj_ct_core_cp_element_group_312 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(312), clk => clk, reset => reset); --
    end block;
    -- CP-element group 313:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	233 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (1) 
      -- CP-element group 313: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_sample_start__ps
      -- 
    ct_core_CP_34_elements(313) <= ct_core_CP_34_elements(233);
    -- CP-element group 314:  join  transition  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	234 
    -- CP-element group 314:  members (1) 
      -- CP-element group 314: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_sample_completed__ps
      -- 
    -- Element group ct_core_CP_34_elements(314) is bound as output of CP function.
    -- CP-element group 315:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	235 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (1) 
      -- CP-element group 315: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_update_start__ps
      -- 
    ct_core_CP_34_elements(315) <= ct_core_CP_34_elements(235);
    -- CP-element group 316:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	236 
    -- CP-element group 316: 	362 
    -- CP-element group 316: marked-successors 
    -- CP-element group 316: 	312 
    -- CP-element group 316:  members (2) 
      -- CP-element group 316: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_update_completed__ps
      -- CP-element group 316: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_update_completed_
      -- 
    -- Element group ct_core_CP_34_elements(316) is bound as output of CP function.
    -- CP-element group 317:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	229 
    -- CP-element group 317: successors 
    -- CP-element group 317:  members (1) 
      -- CP-element group 317: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_loopback_trigger
      -- 
    ct_core_CP_34_elements(317) <= ct_core_CP_34_elements(229);
    -- CP-element group 318:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (2) 
      -- CP-element group 318: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_loopback_sample_req_ps
      -- CP-element group 318: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_loopback_sample_req
      -- 
    phi_stmt_974_loopback_sample_req_2036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_974_loopback_sample_req_2036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(318), ack => phi_stmt_974_req_1); -- 
    -- Element group ct_core_CP_34_elements(318) is bound as output of CP function.
    -- CP-element group 319:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	230 
    -- CP-element group 319: successors 
    -- CP-element group 319:  members (1) 
      -- CP-element group 319: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_entry_trigger
      -- 
    ct_core_CP_34_elements(319) <= ct_core_CP_34_elements(230);
    -- CP-element group 320:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (2) 
      -- CP-element group 320: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_entry_sample_req
      -- CP-element group 320: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_entry_sample_req_ps
      -- 
    phi_stmt_974_entry_sample_req_2039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_974_entry_sample_req_2039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(320), ack => phi_stmt_974_req_0); -- 
    -- Element group ct_core_CP_34_elements(320) is bound as output of CP function.
    -- CP-element group 321:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: successors 
    -- CP-element group 321:  members (2) 
      -- CP-element group 321: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_phi_mux_ack_ps
      -- CP-element group 321: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_974_phi_mux_ack
      -- 
    phi_stmt_974_phi_mux_ack_2042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_974_ack_0, ack => ct_core_CP_34_elements(321)); -- 
    -- CP-element group 322:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (4) 
      -- CP-element group 322: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_Sample/req
      -- CP-element group 322: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_sample_start__ps
      -- 
    req_2055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(322), ack => add_dest_dim1_init_951_976_buf_req_0); -- 
    -- Element group ct_core_CP_34_elements(322) is bound as output of CP function.
    -- CP-element group 323:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (4) 
      -- CP-element group 323: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_Update/req
      -- CP-element group 323: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_update_start_
      -- CP-element group 323: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_update_start__ps
      -- 
    req_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(323), ack => add_dest_dim1_init_951_976_buf_req_1); -- 
    -- Element group ct_core_CP_34_elements(323) is bound as output of CP function.
    -- CP-element group 324:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: successors 
    -- CP-element group 324:  members (4) 
      -- CP-element group 324: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_Sample/ack
      -- CP-element group 324: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_sample_completed_
      -- CP-element group 324: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_sample_completed__ps
      -- 
    ack_2056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim1_init_951_976_buf_ack_0, ack => ct_core_CP_34_elements(324)); -- 
    -- CP-element group 325:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325:  members (4) 
      -- CP-element group 325: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_Update/ack
      -- CP-element group 325: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_update_completed_
      -- CP-element group 325: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_dest_dim1_init_976_update_completed__ps
      -- 
    ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => add_dest_dim1_init_951_976_buf_ack_1, ack => ct_core_CP_34_elements(325)); -- 
    -- CP-element group 326:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (4) 
      -- CP-element group 326: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_Sample/req
      -- CP-element group 326: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_sample_start__ps
      -- 
    req_2073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(326), ack => next_add_dest_dim1_1121_977_buf_req_0); -- 
    -- Element group ct_core_CP_34_elements(326) is bound as output of CP function.
    -- CP-element group 327:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	329 
    -- CP-element group 327:  members (4) 
      -- CP-element group 327: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_Update/req
      -- CP-element group 327: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_update_start_
      -- CP-element group 327: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_update_start__ps
      -- 
    req_2078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(327), ack => next_add_dest_dim1_1121_977_buf_req_1); -- 
    -- Element group ct_core_CP_34_elements(327) is bound as output of CP function.
    -- CP-element group 328:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: successors 
    -- CP-element group 328:  members (4) 
      -- CP-element group 328: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_Sample/ack
      -- CP-element group 328: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_Sample/$exit
      -- CP-element group 328: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_sample_completed_
      -- CP-element group 328: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_sample_completed__ps
      -- 
    ack_2074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim1_1121_977_buf_ack_0, ack => ct_core_CP_34_elements(328)); -- 
    -- CP-element group 329:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	327 
    -- CP-element group 329: successors 
    -- CP-element group 329:  members (4) 
      -- CP-element group 329: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_Update/ack
      -- CP-element group 329: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_Update/$exit
      -- CP-element group 329: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_update_completed_
      -- CP-element group 329: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_dest_dim1_977_update_completed__ps
      -- 
    ack_2079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_dest_dim1_1121_977_buf_ack_1, ack => ct_core_CP_34_elements(329)); -- 
    -- CP-element group 330:  join  transition  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	231 
    -- CP-element group 330: marked-predecessors 
    -- CP-element group 330: 	234 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	233 
    -- CP-element group 330:  members (1) 
      -- CP-element group 330: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_sample_start_
      -- 
    ct_core_cp_element_group_330: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_330"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(234);
      gj_ct_core_cp_element_group_330 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(330), clk => clk, reset => reset); --
    end block;
    -- CP-element group 331:  join  transition  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	231 
    -- CP-element group 331: marked-predecessors 
    -- CP-element group 331: 	335 
    -- CP-element group 331: 	352 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	235 
    -- CP-element group 331:  members (1) 
      -- CP-element group 331: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_update_start_
      -- 
    ct_core_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(335) & ct_core_CP_34_elements(352);
      gj_ct_core_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	233 
    -- CP-element group 332: successors 
    -- CP-element group 332:  members (1) 
      -- CP-element group 332: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_sample_start__ps
      -- 
    ct_core_CP_34_elements(332) <= ct_core_CP_34_elements(233);
    -- CP-element group 333:  join  transition  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	234 
    -- CP-element group 333:  members (1) 
      -- CP-element group 333: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_sample_completed__ps
      -- 
    -- Element group ct_core_CP_34_elements(333) is bound as output of CP function.
    -- CP-element group 334:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	235 
    -- CP-element group 334: successors 
    -- CP-element group 334:  members (1) 
      -- CP-element group 334: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_update_start__ps
      -- 
    ct_core_CP_34_elements(334) <= ct_core_CP_34_elements(235);
    -- CP-element group 335:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	236 
    -- CP-element group 335: 	352 
    -- CP-element group 335: marked-successors 
    -- CP-element group 335: 	331 
    -- CP-element group 335:  members (15) 
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_scale_1/$entry
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_scale_1/scale_rename_ack
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_update_completed_
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_update_completed__ps
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_scale_1/$exit
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_scale_1/scale_rename_req
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_final_index_sum_regn_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_resize_1/index_resize_ack
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_resize_1/index_resize_req
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_resize_1/$exit
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_resize_1/$entry
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_computed_1
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_scaled_1
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_index_resized_1
      -- CP-element group 335: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_final_index_sum_regn_Sample/req
      -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(335), ack => array_obj_ref_1013_index_offset_req_0); -- 
    -- Element group ct_core_CP_34_elements(335) is bound as output of CP function.
    -- CP-element group 336:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	229 
    -- CP-element group 336: successors 
    -- CP-element group 336:  members (1) 
      -- CP-element group 336: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_loopback_trigger
      -- 
    ct_core_CP_34_elements(336) <= ct_core_CP_34_elements(229);
    -- CP-element group 337:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: successors 
    -- CP-element group 337:  members (2) 
      -- CP-element group 337: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_loopback_sample_req
      -- CP-element group 337: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_loopback_sample_req_ps
      -- 
    phi_stmt_978_loopback_sample_req_2090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_978_loopback_sample_req_2090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(337), ack => phi_stmt_978_req_1); -- 
    -- Element group ct_core_CP_34_elements(337) is bound as output of CP function.
    -- CP-element group 338:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	230 
    -- CP-element group 338: successors 
    -- CP-element group 338:  members (1) 
      -- CP-element group 338: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_entry_trigger
      -- 
    ct_core_CP_34_elements(338) <= ct_core_CP_34_elements(230);
    -- CP-element group 339:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: successors 
    -- CP-element group 339:  members (2) 
      -- CP-element group 339: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_entry_sample_req_ps
      -- CP-element group 339: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_entry_sample_req
      -- 
    phi_stmt_978_entry_sample_req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_978_entry_sample_req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(339), ack => phi_stmt_978_req_0); -- 
    -- Element group ct_core_CP_34_elements(339) is bound as output of CP function.
    -- CP-element group 340:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: successors 
    -- CP-element group 340:  members (2) 
      -- CP-element group 340: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_phi_mux_ack_ps
      -- CP-element group 340: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/phi_stmt_978_phi_mux_ack
      -- 
    phi_stmt_978_phi_mux_ack_2096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_978_ack_0, ack => ct_core_CP_34_elements(340)); -- 
    -- CP-element group 341:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: successors 
    -- CP-element group 341:  members (4) 
      -- CP-element group 341: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_src_init_980_sample_completed__ps
      -- CP-element group 341: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_src_init_980_sample_start__ps
      -- CP-element group 341: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_src_init_980_sample_start_
      -- CP-element group 341: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_src_init_980_sample_completed_
      -- 
    -- Element group ct_core_CP_34_elements(341) is bound as output of CP function.
    -- CP-element group 342:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (2) 
      -- CP-element group 342: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_src_init_980_update_start__ps
      -- CP-element group 342: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_src_init_980_update_start_
      -- 
    -- Element group ct_core_CP_34_elements(342) is bound as output of CP function.
    -- CP-element group 343:  join  transition  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	344 
    -- CP-element group 343: successors 
    -- CP-element group 343:  members (1) 
      -- CP-element group 343: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_src_init_980_update_completed__ps
      -- 
    ct_core_CP_34_elements(343) <= ct_core_CP_34_elements(344);
    -- CP-element group 344:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	343 
    -- CP-element group 344:  members (1) 
      -- CP-element group 344: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_add_src_init_980_update_completed_
      -- 
    -- Element group ct_core_CP_34_elements(344) is a control-delay.
    cp_element_344_delay: control_delay_element  generic map(name => " 344_delay", delay_value => 1)  port map(req => ct_core_CP_34_elements(342), ack => ct_core_CP_34_elements(344), clk => clk, reset =>reset);
    -- CP-element group 345:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (4) 
      -- CP-element group 345: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_Sample/req
      -- CP-element group 345: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_sample_start_
      -- CP-element group 345: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_sample_start__ps
      -- 
    req_2117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(345), ack => next_add_src_1111_981_buf_req_0); -- 
    -- Element group ct_core_CP_34_elements(345) is bound as output of CP function.
    -- CP-element group 346:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (4) 
      -- CP-element group 346: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_Update/$entry
      -- CP-element group 346: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_Update/req
      -- CP-element group 346: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_update_start_
      -- CP-element group 346: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_update_start__ps
      -- 
    req_2122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(346), ack => next_add_src_1111_981_buf_req_1); -- 
    -- Element group ct_core_CP_34_elements(346) is bound as output of CP function.
    -- CP-element group 347:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347:  members (4) 
      -- CP-element group 347: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_sample_completed__ps
      -- 
    ack_2118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_src_1111_981_buf_ack_0, ack => ct_core_CP_34_elements(347)); -- 
    -- CP-element group 348:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: successors 
    -- CP-element group 348:  members (4) 
      -- CP-element group 348: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_Update/ack
      -- CP-element group 348: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/R_next_add_src_981_update_completed__ps
      -- 
    ack_2123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_src_1111_981_buf_ack_1, ack => ct_core_CP_34_elements(348)); -- 
    -- CP-element group 349:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	353 
    -- CP-element group 349: marked-predecessors 
    -- CP-element group 349: 	354 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	354 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_request/$entry
      -- CP-element group 349: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_sample_start_
      -- CP-element group 349: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_request/req
      -- 
    req_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(349), ack => addr_of_1014_final_reg_req_0); -- 
    ct_core_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(353) & ct_core_CP_34_elements(354);
      gj_ct_core_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	231 
    -- CP-element group 350: marked-predecessors 
    -- CP-element group 350: 	358 
    -- CP-element group 350: 	355 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	355 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_update_start_
      -- CP-element group 350: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_complete/req
      -- CP-element group 350: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_complete/$entry
      -- 
    req_2169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(350), ack => addr_of_1014_final_reg_req_1); -- 
    ct_core_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(358) & ct_core_CP_34_elements(355);
      gj_ct_core_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	231 
    -- CP-element group 351: marked-predecessors 
    -- CP-element group 351: 	353 
    -- CP-element group 351: 	354 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_final_index_sum_regn_update_start
      -- CP-element group 351: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_final_index_sum_regn_Update/req
      -- CP-element group 351: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_final_index_sum_regn_Update/$entry
      -- 
    req_2154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(351), ack => array_obj_ref_1013_index_offset_req_1); -- 
    ct_core_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(353) & ct_core_CP_34_elements(354);
      gj_ct_core_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	335 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	393 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	331 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_final_index_sum_regn_sample_complete
      -- CP-element group 352: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_final_index_sum_regn_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_final_index_sum_regn_Sample/$exit
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1013_index_offset_ack_0, ack => ct_core_CP_34_elements(352)); -- 
    -- CP-element group 353:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	349 
    -- CP-element group 353: marked-successors 
    -- CP-element group 353: 	351 
    -- CP-element group 353:  members (8) 
      -- CP-element group 353: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_base_plus_offset/sum_rename_ack
      -- CP-element group 353: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_base_plus_offset/$entry
      -- CP-element group 353: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_base_plus_offset/sum_rename_req
      -- CP-element group 353: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_base_plus_offset/$exit
      -- CP-element group 353: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_final_index_sum_regn_Update/ack
      -- CP-element group 353: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_offset_calculated
      -- CP-element group 353: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_root_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1013_final_index_sum_regn_Update/$exit
      -- 
    ack_2155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1013_index_offset_ack_1, ack => ct_core_CP_34_elements(353)); -- 
    -- CP-element group 354:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	349 
    -- CP-element group 354: successors 
    -- CP-element group 354: marked-successors 
    -- CP-element group 354: 	349 
    -- CP-element group 354: 	351 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_request/$exit
      -- CP-element group 354: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_request/ack
      -- 
    ack_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1014_final_reg_ack_0, ack => ct_core_CP_34_elements(354)); -- 
    -- CP-element group 355:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	350 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355: marked-successors 
    -- CP-element group 355: 	350 
    -- CP-element group 355:  members (19) 
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_base_plus_offset/$entry
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_base_addr_resize/base_resize_req
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_base_addr_resize/base_resize_ack
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_base_addr_resize/$exit
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_base_addr_resize/$entry
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_base_address_resized
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_root_address_calculated
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_word_address_calculated
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_base_address_calculated
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_word_addrgen/root_register_ack
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_complete/ack
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_word_addrgen/root_register_req
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_word_addrgen/$exit
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_word_addrgen/$entry
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1014_complete/$exit
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_base_plus_offset/sum_rename_ack
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_base_plus_offset/sum_rename_req
      -- CP-element group 355: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_base_plus_offset/$exit
      -- 
    ack_2170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1014_final_reg_ack_1, ack => ct_core_CP_34_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: marked-predecessors 
    -- CP-element group 356: 	358 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	358 
    -- CP-element group 356:  members (5) 
      -- CP-element group 356: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Sample/word_access_start/word_0/rr
      -- CP-element group 356: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Sample/word_access_start/word_0/$entry
      -- CP-element group 356: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Sample/word_access_start/$entry
      -- CP-element group 356: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_sample_start_
      -- 
    rr_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(356), ack => ptr_deref_1018_load_0_req_0); -- 
    ct_core_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(355) & ct_core_CP_34_elements(358);
      gj_ct_core_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: marked-predecessors 
    -- CP-element group 357: 	374 
    -- CP-element group 357: 	359 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (5) 
      -- CP-element group 357: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/word_access_complete/$entry
      -- CP-element group 357: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_update_start_
      -- CP-element group 357: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/word_access_complete/word_0/cr
      -- CP-element group 357: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/word_access_complete/word_0/$entry
      -- 
    cr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(357), ack => ptr_deref_1018_load_0_req_1); -- 
    ct_core_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(374) & ct_core_CP_34_elements(359);
      gj_ct_core_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	356 
    -- CP-element group 358: successors 
    -- CP-element group 358: marked-successors 
    -- CP-element group 358: 	350 
    -- CP-element group 358: 	356 
    -- CP-element group 358:  members (5) 
      -- CP-element group 358: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Sample/word_access_start/word_0/ra
      -- CP-element group 358: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Sample/word_access_start/word_0/$exit
      -- CP-element group 358: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Sample/word_access_start/$exit
      -- CP-element group 358: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Sample/$exit
      -- CP-element group 358: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_sample_completed_
      -- 
    ra_2204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1018_load_0_ack_0, ack => ct_core_CP_34_elements(358)); -- 
    -- CP-element group 359:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	372 
    -- CP-element group 359: marked-successors 
    -- CP-element group 359: 	357 
    -- CP-element group 359:  members (9) 
      -- CP-element group 359: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/$exit
      -- CP-element group 359: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/word_access_complete/$exit
      -- CP-element group 359: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/ptr_deref_1018_Merge/merge_ack
      -- CP-element group 359: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_update_completed_
      -- CP-element group 359: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/ptr_deref_1018_Merge/merge_req
      -- CP-element group 359: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/ptr_deref_1018_Merge/$exit
      -- CP-element group 359: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/ptr_deref_1018_Merge/$entry
      -- CP-element group 359: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/word_access_complete/word_0/ca
      -- CP-element group 359: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1018_Update/word_access_complete/word_0/$exit
      -- 
    ca_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1018_load_0_ack_1, ack => ct_core_CP_34_elements(359)); -- 
    -- CP-element group 360:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	365 
    -- CP-element group 360: marked-predecessors 
    -- CP-element group 360: 	366 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	366 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_request/req
      -- CP-element group 360: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_request/$entry
      -- 
    req_2260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(360), ack => addr_of_1026_final_reg_req_0); -- 
    ct_core_cp_element_group_360: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_360"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(365) & ct_core_CP_34_elements(366);
      gj_ct_core_cp_element_group_360 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(360), clk => clk, reset => reset); --
    end block;
    -- CP-element group 361:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	231 
    -- CP-element group 361: marked-predecessors 
    -- CP-element group 361: 	367 
    -- CP-element group 361: 	370 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	367 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_complete/req
      -- CP-element group 361: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_complete/$entry
      -- CP-element group 361: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_update_start_
      -- 
    req_2265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(361), ack => addr_of_1026_final_reg_req_1); -- 
    ct_core_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(367) & ct_core_CP_34_elements(370);
      gj_ct_core_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	278 
    -- CP-element group 362: 	297 
    -- CP-element group 362: 	316 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (13) 
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_final_index_sum_regn_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_resized_1
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_scale_1/scale_rename_ack
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_scale_1/scale_rename_req
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_scale_1/$exit
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_scale_1/$entry
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_resize_1/index_resize_ack
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_resize_1/index_resize_req
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_resize_1/$exit
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_resize_1/$entry
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_final_index_sum_regn_Sample/req
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_computed_1
      -- CP-element group 362: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_index_scaled_1
      -- 
    req_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(362), ack => array_obj_ref_1025_index_offset_req_0); -- 
    ct_core_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(278) & ct_core_CP_34_elements(297) & ct_core_CP_34_elements(316);
      gj_ct_core_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	231 
    -- CP-element group 363: marked-predecessors 
    -- CP-element group 363: 	365 
    -- CP-element group 363: 	366 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	365 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_final_index_sum_regn_update_start
      -- CP-element group 363: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_final_index_sum_regn_Update/req
      -- CP-element group 363: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_final_index_sum_regn_Update/$entry
      -- 
    req_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(363), ack => array_obj_ref_1025_index_offset_req_1); -- 
    ct_core_cp_element_group_363: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_363"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(365) & ct_core_CP_34_elements(366);
      gj_ct_core_cp_element_group_363 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 364:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	393 
    -- CP-element group 364: marked-successors 
    -- CP-element group 364: 	274 
    -- CP-element group 364: 	293 
    -- CP-element group 364: 	312 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_final_index_sum_regn_sample_complete
      -- CP-element group 364: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_final_index_sum_regn_Sample/ack
      -- CP-element group 364: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_final_index_sum_regn_Sample/$exit
      -- 
    ack_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1025_index_offset_ack_0, ack => ct_core_CP_34_elements(364)); -- 
    -- CP-element group 365:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	363 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	360 
    -- CP-element group 365: marked-successors 
    -- CP-element group 365: 	363 
    -- CP-element group 365:  members (8) 
      -- CP-element group 365: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_base_plus_offset/$entry
      -- CP-element group 365: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_root_address_calculated
      -- CP-element group 365: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_base_plus_offset/sum_rename_ack
      -- CP-element group 365: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_base_plus_offset/sum_rename_req
      -- CP-element group 365: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_base_plus_offset/$exit
      -- CP-element group 365: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_offset_calculated
      -- CP-element group 365: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_final_index_sum_regn_Update/ack
      -- CP-element group 365: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/array_obj_ref_1025_final_index_sum_regn_Update/$exit
      -- 
    ack_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1025_index_offset_ack_1, ack => ct_core_CP_34_elements(365)); -- 
    -- CP-element group 366:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	360 
    -- CP-element group 366: successors 
    -- CP-element group 366: marked-successors 
    -- CP-element group 366: 	360 
    -- CP-element group 366: 	363 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_request/ack
      -- CP-element group 366: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_sample_completed_
      -- CP-element group 366: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_request/$exit
      -- 
    ack_2261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1026_final_reg_ack_0, ack => ct_core_CP_34_elements(366)); -- 
    -- CP-element group 367:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	361 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367: marked-successors 
    -- CP-element group 367: 	361 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_complete/ack
      -- CP-element group 367: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_complete/$exit
      -- CP-element group 367: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/addr_of_1026_update_completed_
      -- 
    ack_2266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1026_final_reg_ack_1, ack => ct_core_CP_34_elements(367)); -- 
    -- CP-element group 368:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: marked-predecessors 
    -- CP-element group 368: 	370 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	370 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_Sample/$entry
      -- CP-element group 368: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_Sample/req
      -- CP-element group 368: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_sample_start_
      -- 
    req_2274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(368), ack => W_ov_1028_delayed_6_0_1028_inst_req_0); -- 
    ct_core_cp_element_group_368: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_368"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(367) & ct_core_CP_34_elements(370);
      gj_ct_core_cp_element_group_368 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 369:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: marked-predecessors 
    -- CP-element group 369: 	371 
    -- CP-element group 369: 	374 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	371 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_Update/req
      -- CP-element group 369: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_Update/$entry
      -- CP-element group 369: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_update_start_
      -- 
    req_2279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(369), ack => W_ov_1028_delayed_6_0_1028_inst_req_1); -- 
    ct_core_cp_element_group_369: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_369"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(371) & ct_core_CP_34_elements(374);
      gj_ct_core_cp_element_group_369 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(369), clk => clk, reset => reset); --
    end block;
    -- CP-element group 370:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	368 
    -- CP-element group 370: successors 
    -- CP-element group 370: marked-successors 
    -- CP-element group 370: 	361 
    -- CP-element group 370: 	368 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_Sample/ack
      -- CP-element group 370: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_sample_completed_
      -- 
    ack_2275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ov_1028_delayed_6_0_1028_inst_ack_0, ack => ct_core_CP_34_elements(370)); -- 
    -- CP-element group 371:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	369 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371: marked-successors 
    -- CP-element group 371: 	369 
    -- CP-element group 371:  members (19) 
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_Update/ack
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1030_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_base_address_calculated
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_word_address_calculated
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_root_address_calculated
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_base_address_resized
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_base_addr_resize/$entry
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_base_addr_resize/$exit
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_base_addr_resize/base_resize_req
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_base_addr_resize/base_resize_ack
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_base_plus_offset/$entry
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_base_plus_offset/$exit
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_base_plus_offset/sum_rename_req
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_base_plus_offset/sum_rename_ack
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_word_addrgen/$entry
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_word_addrgen/$exit
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_word_addrgen/root_register_req
      -- CP-element group 371: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_word_addrgen/root_register_ack
      -- 
    ack_2280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ov_1028_delayed_6_0_1028_inst_ack_1, ack => ct_core_CP_34_elements(371)); -- 
    -- CP-element group 372:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: 	359 
    -- CP-element group 372: marked-predecessors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372:  members (9) 
      -- CP-element group 372: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_sample_start_
      -- CP-element group 372: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/ptr_deref_1032_Split/$entry
      -- CP-element group 372: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/ptr_deref_1032_Split/$exit
      -- CP-element group 372: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/ptr_deref_1032_Split/split_req
      -- CP-element group 372: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/ptr_deref_1032_Split/split_ack
      -- CP-element group 372: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/word_access_start/$entry
      -- CP-element group 372: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/word_access_start/word_0/$entry
      -- CP-element group 372: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/word_access_start/word_0/rr
      -- 
    rr_2318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(372), ack => ptr_deref_1032_store_0_req_0); -- 
    ct_core_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(371) & ct_core_CP_34_elements(359) & ct_core_CP_34_elements(374);
      gj_ct_core_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: marked-predecessors 
    -- CP-element group 373: 	375 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (5) 
      -- CP-element group 373: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_update_start_
      -- CP-element group 373: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Update/word_access_complete/$entry
      -- CP-element group 373: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Update/word_access_complete/word_0/$entry
      -- CP-element group 373: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Update/word_access_complete/word_0/cr
      -- 
    cr_2329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(373), ack => ptr_deref_1032_store_0_req_1); -- 
    ct_core_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ct_core_CP_34_elements(375);
      gj_ct_core_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: marked-successors 
    -- CP-element group 374: 	369 
    -- CP-element group 374: 	372 
    -- CP-element group 374: 	357 
    -- CP-element group 374:  members (5) 
      -- CP-element group 374: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/$exit
      -- CP-element group 374: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/word_access_start/$exit
      -- CP-element group 374: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/word_access_start/word_0/$exit
      -- CP-element group 374: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Sample/word_access_start/word_0/ra
      -- 
    ra_2319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1032_store_0_ack_0, ack => ct_core_CP_34_elements(374)); -- 
    -- CP-element group 375:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	393 
    -- CP-element group 375: marked-successors 
    -- CP-element group 375: 	373 
    -- CP-element group 375:  members (5) 
      -- CP-element group 375: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Update/word_access_complete/$exit
      -- CP-element group 375: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Update/word_access_complete/word_0/$exit
      -- CP-element group 375: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/ptr_deref_1032_Update/word_access_complete/word_0/ca
      -- 
    ca_2330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1032_store_0_ack_1, ack => ct_core_CP_34_elements(375)); -- 
    -- CP-element group 376:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	231 
    -- CP-element group 376: marked-predecessors 
    -- CP-element group 376: 	378 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	378 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_sample_start_
      -- CP-element group 376: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_Sample/req
      -- 
    req_2338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(376), ack => W_dim2_limit_1039_delayed_1_0_1040_inst_req_0); -- 
    ct_core_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(378);
      gj_ct_core_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	234 
    -- CP-element group 377: marked-predecessors 
    -- CP-element group 377: 	379 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_update_start_
      -- CP-element group 377: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_Update/$entry
      -- CP-element group 377: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_Update/req
      -- 
    req_2343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(377), ack => W_dim2_limit_1039_delayed_1_0_1040_inst_req_1); -- 
    ct_core_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(234) & ct_core_CP_34_elements(379);
      gj_ct_core_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	376 
    -- CP-element group 378: successors 
    -- CP-element group 378: marked-successors 
    -- CP-element group 378: 	376 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_Sample/ack
      -- 
    ack_2339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dim2_limit_1039_delayed_1_0_1040_inst_ack_0, ack => ct_core_CP_34_elements(378)); -- 
    -- CP-element group 379:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	232 
    -- CP-element group 379: marked-successors 
    -- CP-element group 379: 	237 
    -- CP-element group 379: 	254 
    -- CP-element group 379: 	273 
    -- CP-element group 379: 	292 
    -- CP-element group 379: 	311 
    -- CP-element group 379: 	377 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1042_Update/ack
      -- 
    ack_2344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dim2_limit_1039_delayed_1_0_1040_inst_ack_1, ack => ct_core_CP_34_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	231 
    -- CP-element group 380: marked-predecessors 
    -- CP-element group 380: 	382 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_sample_start_
      -- CP-element group 380: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_Sample/$entry
      -- CP-element group 380: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_Sample/rr
      -- 
    rr_2352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(380), ack => SUB_u16_u16_1051_inst_req_0); -- 
    ct_core_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(382);
      gj_ct_core_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	234 
    -- CP-element group 381: marked-predecessors 
    -- CP-element group 381: 	383 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	383 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_update_start_
      -- CP-element group 381: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_Update/$entry
      -- CP-element group 381: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_Update/cr
      -- 
    cr_2357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(381), ack => SUB_u16_u16_1051_inst_req_1); -- 
    ct_core_cp_element_group_381: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_381"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(234) & ct_core_CP_34_elements(383);
      gj_ct_core_cp_element_group_381 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(381), clk => clk, reset => reset); --
    end block;
    -- CP-element group 382:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382: marked-successors 
    -- CP-element group 382: 	380 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_Sample/ra
      -- 
    ra_2353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1051_inst_ack_0, ack => ct_core_CP_34_elements(382)); -- 
    -- CP-element group 383:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	381 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	232 
    -- CP-element group 383: marked-successors 
    -- CP-element group 383: 	237 
    -- CP-element group 383: 	254 
    -- CP-element group 383: 	292 
    -- CP-element group 383: 	311 
    -- CP-element group 383: 	381 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1051_Update/ca
      -- 
    ca_2358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1051_inst_ack_1, ack => ct_core_CP_34_elements(383)); -- 
    -- CP-element group 384:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	231 
    -- CP-element group 384: marked-predecessors 
    -- CP-element group 384: 	386 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	386 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_sample_start_
      -- CP-element group 384: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_Sample/$entry
      -- CP-element group 384: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_Sample/req
      -- 
    req_2366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(384), ack => W_nid1_true3_1092_delayed_1_0_1099_inst_req_0); -- 
    ct_core_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(386);
      gj_ct_core_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	234 
    -- CP-element group 385: marked-predecessors 
    -- CP-element group 385: 	387 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	387 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_update_start_
      -- CP-element group 385: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_Update/$entry
      -- CP-element group 385: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_Update/req
      -- 
    req_2371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(385), ack => W_nid1_true3_1092_delayed_1_0_1099_inst_req_1); -- 
    ct_core_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(234) & ct_core_CP_34_elements(387);
      gj_ct_core_cp_element_group_385 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	384 
    -- CP-element group 386: successors 
    -- CP-element group 386: marked-successors 
    -- CP-element group 386: 	384 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_Sample/ack
      -- 
    ack_2367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_nid1_true3_1092_delayed_1_0_1099_inst_ack_0, ack => ct_core_CP_34_elements(386)); -- 
    -- CP-element group 387:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	385 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	393 
    -- CP-element group 387: marked-successors 
    -- CP-element group 387: 	311 
    -- CP-element group 387: 	385 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/assign_stmt_1101_Update/ack
      -- 
    ack_2372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_nid1_true3_1092_delayed_1_0_1099_inst_ack_1, ack => ct_core_CP_34_elements(387)); -- 
    -- CP-element group 388:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	231 
    -- CP-element group 388: marked-predecessors 
    -- CP-element group 388: 	390 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	390 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_sample_start_
      -- CP-element group 388: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_Sample/$entry
      -- CP-element group 388: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_Sample/rr
      -- 
    rr_2380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(388), ack => SUB_u16_u16_1153_inst_req_0); -- 
    ct_core_cp_element_group_388: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_388"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(231) & ct_core_CP_34_elements(390);
      gj_ct_core_cp_element_group_388 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(388), clk => clk, reset => reset); --
    end block;
    -- CP-element group 389:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: marked-predecessors 
    -- CP-element group 389: 	391 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	391 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_update_start_
      -- CP-element group 389: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_Update/$entry
      -- CP-element group 389: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_Update/cr
      -- 
    cr_2385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(389), ack => SUB_u16_u16_1153_inst_req_1); -- 
    ct_core_cp_element_group_389: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_389"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ct_core_CP_34_elements(391);
      gj_ct_core_cp_element_group_389 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(389), clk => clk, reset => reset); --
    end block;
    -- CP-element group 390:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	388 
    -- CP-element group 390: successors 
    -- CP-element group 390: marked-successors 
    -- CP-element group 390: 	388 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_Sample/ra
      -- 
    ra_2381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1153_inst_ack_0, ack => ct_core_CP_34_elements(390)); -- 
    -- CP-element group 391:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	389 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	232 
    -- CP-element group 391: marked-successors 
    -- CP-element group 391: 	389 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/SUB_u16_u16_1153_Update/ca
      -- 
    ca_2386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1153_inst_ack_1, ack => ct_core_CP_34_elements(391)); -- 
    -- CP-element group 392:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	231 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	232 
    -- CP-element group 392:  members (1) 
      -- CP-element group 392: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group ct_core_CP_34_elements(392) is a control-delay.
    cp_element_392_delay: control_delay_element  generic map(name => " 392_delay", delay_value => 1)  port map(req => ct_core_CP_34_elements(231), ack => ct_core_CP_34_elements(392), clk => clk, reset =>reset);
    -- CP-element group 393:  join  transition  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	234 
    -- CP-element group 393: 	364 
    -- CP-element group 393: 	375 
    -- CP-element group 393: 	387 
    -- CP-element group 393: 	352 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	228 
    -- CP-element group 393:  members (1) 
      -- CP-element group 393: 	 branch_block_stmt_25/do_while_stmt_956/do_while_stmt_956_loop_body/$exit
      -- 
    ct_core_cp_element_group_393: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_393"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(234) & ct_core_CP_34_elements(364) & ct_core_CP_34_elements(375) & ct_core_CP_34_elements(387) & ct_core_CP_34_elements(352);
      gj_ct_core_cp_element_group_393 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(393), clk => clk, reset => reset); --
    end block;
    -- CP-element group 394:  transition  input  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	227 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (2) 
      -- CP-element group 394: 	 branch_block_stmt_25/do_while_stmt_956/loop_exit/$exit
      -- CP-element group 394: 	 branch_block_stmt_25/do_while_stmt_956/loop_exit/ack
      -- 
    ack_2391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_956_branch_ack_0, ack => ct_core_CP_34_elements(394)); -- 
    -- CP-element group 395:  transition  input  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	227 
    -- CP-element group 395: successors 
    -- CP-element group 395:  members (2) 
      -- CP-element group 395: 	 branch_block_stmt_25/do_while_stmt_956/loop_taken/$exit
      -- CP-element group 395: 	 branch_block_stmt_25/do_while_stmt_956/loop_taken/ack
      -- 
    ack_2395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_956_branch_ack_1, ack => ct_core_CP_34_elements(395)); -- 
    -- CP-element group 396:  transition  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	225 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	1 
    -- CP-element group 396:  members (1) 
      -- CP-element group 396: 	 branch_block_stmt_25/do_while_stmt_956/$exit
      -- 
    ct_core_CP_34_elements(396) <= ct_core_CP_34_elements(225);
    -- CP-element group 397:  transition  input  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	1 
    -- CP-element group 397: successors 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_sample_completed_
      -- CP-element group 397: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_Sample/$exit
      -- CP-element group 397: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_Sample/cra
      -- 
    cra_2408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1170_call_ack_0, ack => ct_core_CP_34_elements(397)); -- 
    -- CP-element group 398:  transition  input  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	1 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	401 
    -- CP-element group 398:  members (6) 
      -- CP-element group 398: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_update_completed_
      -- CP-element group 398: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_Update/$exit
      -- CP-element group 398: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/call_stmt_1170_Update/cca
      -- CP-element group 398: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_Sample/rr
      -- 
    cca_2413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1170_call_ack_1, ack => ct_core_CP_34_elements(398)); -- 
    rr_2435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(398), ack => type_cast_1180_inst_req_0); -- 
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	1 
    -- CP-element group 399: successors 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_sample_completed_
      -- CP-element group 399: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_Sample/$exit
      -- CP-element group 399: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_Sample/ra
      -- 
    ra_2422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1175_inst_ack_0, ack => ct_core_CP_34_elements(399)); -- 
    -- CP-element group 400:  transition  input  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	1 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	403 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_update_completed_
      -- CP-element group 400: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_Update/$exit
      -- CP-element group 400: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1175_Update/ca
      -- 
    ca_2427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1175_inst_ack_1, ack => ct_core_CP_34_elements(400)); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	398 
    -- CP-element group 401: successors 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_sample_completed_
      -- CP-element group 401: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_Sample/$exit
      -- CP-element group 401: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_Sample/ra
      -- 
    ra_2436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1180_inst_ack_0, ack => ct_core_CP_34_elements(401)); -- 
    -- CP-element group 402:  transition  input  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	1 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_update_completed_
      -- CP-element group 402: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_Update/$exit
      -- CP-element group 402: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/type_cast_1180_Update/ca
      -- 
    ca_2441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1180_inst_ack_1, ack => ct_core_CP_34_elements(402)); -- 
    -- CP-element group 403:  join  fork  transition  place  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	400 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	405 
    -- CP-element group 403: 	406 
    -- CP-element group 403: 	407 
    -- CP-element group 403: 	408 
    -- CP-element group 403: 	409 
    -- CP-element group 403: 	410 
    -- CP-element group 403: 	411 
    -- CP-element group 403: 	412 
    -- CP-element group 403: 	413 
    -- CP-element group 403: 	414 
    -- CP-element group 403: 	415 
    -- CP-element group 403: 	416 
    -- CP-element group 403: 	417 
    -- CP-element group 403: 	418 
    -- CP-element group 403: 	419 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (52) 
      -- CP-element group 403: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186__exit__
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285__entry__
      -- CP-element group 403: 	 branch_block_stmt_25/call_stmt_1170_to_assign_stmt_1186/$exit
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_update_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_Sample/rr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_Update/cr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_update_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_Sample/rr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_Update/cr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_update_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_Sample/rr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_Update/cr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_update_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_Sample/rr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_Update/cr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_update_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_Sample/rr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_Update/cr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_update_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_Sample/rr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_Update/cr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_update_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_Sample/rr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_Update/cr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_update_start_
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_Sample/rr
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_Update/cr
      -- 
    rr_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1190_inst_req_0); -- 
    cr_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1190_inst_req_1); -- 
    rr_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1200_inst_req_0); -- 
    cr_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1200_inst_req_1); -- 
    rr_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1210_inst_req_0); -- 
    cr_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1210_inst_req_1); -- 
    rr_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1220_inst_req_0); -- 
    cr_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1220_inst_req_1); -- 
    rr_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1230_inst_req_0); -- 
    cr_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1230_inst_req_1); -- 
    rr_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1240_inst_req_0); -- 
    cr_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1240_inst_req_1); -- 
    rr_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1250_inst_req_0); -- 
    cr_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1250_inst_req_1); -- 
    rr_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1260_inst_req_0); -- 
    cr_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(403), ack => type_cast_1260_inst_req_1); -- 
    ct_core_cp_element_group_403: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_403"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(400) & ct_core_CP_34_elements(402);
      gj_ct_core_cp_element_group_403 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(403), clk => clk, reset => reset); --
    end block;
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_sample_completed_
      -- CP-element group 404: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_Sample/$exit
      -- CP-element group 404: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_Sample/ra
      -- 
    ra_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1190_inst_ack_0, ack => ct_core_CP_34_elements(404)); -- 
    -- CP-element group 405:  transition  input  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	403 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	440 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_update_completed_
      -- CP-element group 405: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_Update/$exit
      -- CP-element group 405: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1190_Update/ca
      -- 
    ca_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1190_inst_ack_1, ack => ct_core_CP_34_elements(405)); -- 
    -- CP-element group 406:  transition  input  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	403 
    -- CP-element group 406: successors 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_sample_completed_
      -- CP-element group 406: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_Sample/$exit
      -- CP-element group 406: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_Sample/ra
      -- 
    ra_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1200_inst_ack_0, ack => ct_core_CP_34_elements(406)); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	403 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	437 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_update_completed_
      -- CP-element group 407: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_Update/$exit
      -- CP-element group 407: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1200_Update/ca
      -- 
    ca_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1200_inst_ack_1, ack => ct_core_CP_34_elements(407)); -- 
    -- CP-element group 408:  transition  input  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	403 
    -- CP-element group 408: successors 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_sample_completed_
      -- CP-element group 408: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_Sample/$exit
      -- CP-element group 408: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_Sample/ra
      -- 
    ra_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1210_inst_ack_0, ack => ct_core_CP_34_elements(408)); -- 
    -- CP-element group 409:  transition  input  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	403 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	434 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_update_completed_
      -- CP-element group 409: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_Update/$exit
      -- CP-element group 409: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1210_Update/ca
      -- 
    ca_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1210_inst_ack_1, ack => ct_core_CP_34_elements(409)); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	403 
    -- CP-element group 410: successors 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_sample_completed_
      -- CP-element group 410: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_Sample/$exit
      -- CP-element group 410: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_Sample/ra
      -- 
    ra_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_0, ack => ct_core_CP_34_elements(410)); -- 
    -- CP-element group 411:  transition  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	403 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	431 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_update_completed_
      -- CP-element group 411: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_Update/$exit
      -- CP-element group 411: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1220_Update/ca
      -- 
    ca_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_1, ack => ct_core_CP_34_elements(411)); -- 
    -- CP-element group 412:  transition  input  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	403 
    -- CP-element group 412: successors 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_sample_completed_
      -- CP-element group 412: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_Sample/ra
      -- 
    ra_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1230_inst_ack_0, ack => ct_core_CP_34_elements(412)); -- 
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	403 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	428 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_update_completed_
      -- CP-element group 413: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1230_Update/ca
      -- 
    ca_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1230_inst_ack_1, ack => ct_core_CP_34_elements(413)); -- 
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	403 
    -- CP-element group 414: successors 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_sample_completed_
      -- CP-element group 414: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_Sample/$exit
      -- CP-element group 414: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_Sample/ra
      -- 
    ra_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1240_inst_ack_0, ack => ct_core_CP_34_elements(414)); -- 
    -- CP-element group 415:  transition  input  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	403 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	425 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_update_completed_
      -- CP-element group 415: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_Update/$exit
      -- CP-element group 415: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1240_Update/ca
      -- 
    ca_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1240_inst_ack_1, ack => ct_core_CP_34_elements(415)); -- 
    -- CP-element group 416:  transition  input  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	403 
    -- CP-element group 416: successors 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_sample_completed_
      -- CP-element group 416: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_Sample/ra
      -- 
    ra_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1250_inst_ack_0, ack => ct_core_CP_34_elements(416)); -- 
    -- CP-element group 417:  transition  input  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	403 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	422 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_update_completed_
      -- CP-element group 417: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1250_Update/ca
      -- 
    ca_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1250_inst_ack_1, ack => ct_core_CP_34_elements(417)); -- 
    -- CP-element group 418:  transition  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	403 
    -- CP-element group 418: successors 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_sample_completed_
      -- CP-element group 418: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_Sample/$exit
      -- CP-element group 418: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_Sample/ra
      -- 
    ra_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1260_inst_ack_0, ack => ct_core_CP_34_elements(418)); -- 
    -- CP-element group 419:  transition  input  output  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	403 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	420 
    -- CP-element group 419:  members (6) 
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_update_completed_
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_Update/$exit
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/type_cast_1260_Update/ca
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_sample_start_
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_Sample/$entry
      -- CP-element group 419: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_Sample/req
      -- 
    ca_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1260_inst_ack_1, ack => ct_core_CP_34_elements(419)); -- 
    req_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(419), ack => WPIPE_ConvTranspose_output_pipe_1262_inst_req_0); -- 
    -- CP-element group 420:  transition  input  output  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	419 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420:  members (6) 
      -- CP-element group 420: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_sample_completed_
      -- CP-element group 420: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_update_start_
      -- CP-element group 420: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_Sample/$exit
      -- CP-element group 420: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_Sample/ack
      -- CP-element group 420: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_Update/$entry
      -- CP-element group 420: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_Update/req
      -- 
    ack_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1262_inst_ack_0, ack => ct_core_CP_34_elements(420)); -- 
    req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(420), ack => WPIPE_ConvTranspose_output_pipe_1262_inst_req_1); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_update_completed_
      -- CP-element group 421: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_Update/$exit
      -- CP-element group 421: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1262_Update/ack
      -- 
    ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1262_inst_ack_1, ack => ct_core_CP_34_elements(421)); -- 
    -- CP-element group 422:  join  transition  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	417 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_sample_start_
      -- CP-element group 422: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_Sample/$entry
      -- CP-element group 422: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_Sample/req
      -- 
    req_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(422), ack => WPIPE_ConvTranspose_output_pipe_1265_inst_req_0); -- 
    ct_core_cp_element_group_422: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_422"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(417) & ct_core_CP_34_elements(421);
      gj_ct_core_cp_element_group_422 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(422), clk => clk, reset => reset); --
    end block;
    -- CP-element group 423:  transition  input  output  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (6) 
      -- CP-element group 423: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_sample_completed_
      -- CP-element group 423: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_update_start_
      -- CP-element group 423: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_Sample/$exit
      -- CP-element group 423: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_Sample/ack
      -- CP-element group 423: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_Update/$entry
      -- CP-element group 423: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_Update/req
      -- 
    ack_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1265_inst_ack_0, ack => ct_core_CP_34_elements(423)); -- 
    req_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(423), ack => WPIPE_ConvTranspose_output_pipe_1265_inst_req_1); -- 
    -- CP-element group 424:  transition  input  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_update_completed_
      -- CP-element group 424: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_Update/$exit
      -- CP-element group 424: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1265_Update/ack
      -- 
    ack_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1265_inst_ack_1, ack => ct_core_CP_34_elements(424)); -- 
    -- CP-element group 425:  join  transition  output  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	415 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_sample_start_
      -- CP-element group 425: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_Sample/$entry
      -- CP-element group 425: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_Sample/req
      -- 
    req_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(425), ack => WPIPE_ConvTranspose_output_pipe_1268_inst_req_0); -- 
    ct_core_cp_element_group_425: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_425"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(415) & ct_core_CP_34_elements(424);
      gj_ct_core_cp_element_group_425 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(425), clk => clk, reset => reset); --
    end block;
    -- CP-element group 426:  transition  input  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426:  members (6) 
      -- CP-element group 426: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_sample_completed_
      -- CP-element group 426: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_update_start_
      -- CP-element group 426: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_Sample/$exit
      -- CP-element group 426: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_Sample/ack
      -- CP-element group 426: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_Update/$entry
      -- CP-element group 426: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_Update/req
      -- 
    ack_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1268_inst_ack_0, ack => ct_core_CP_34_elements(426)); -- 
    req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(426), ack => WPIPE_ConvTranspose_output_pipe_1268_inst_req_1); -- 
    -- CP-element group 427:  transition  input  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_update_completed_
      -- CP-element group 427: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_Update/$exit
      -- CP-element group 427: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1268_Update/ack
      -- 
    ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1268_inst_ack_1, ack => ct_core_CP_34_elements(427)); -- 
    -- CP-element group 428:  join  transition  output  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	413 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_sample_start_
      -- CP-element group 428: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_Sample/$entry
      -- CP-element group 428: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_Sample/req
      -- 
    req_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(428), ack => WPIPE_ConvTranspose_output_pipe_1271_inst_req_0); -- 
    ct_core_cp_element_group_428: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_428"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(413) & ct_core_CP_34_elements(427);
      gj_ct_core_cp_element_group_428 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(428), clk => clk, reset => reset); --
    end block;
    -- CP-element group 429:  transition  input  output  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	428 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429:  members (6) 
      -- CP-element group 429: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_sample_completed_
      -- CP-element group 429: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_update_start_
      -- CP-element group 429: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_Sample/$exit
      -- CP-element group 429: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_Sample/ack
      -- CP-element group 429: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_Update/$entry
      -- CP-element group 429: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_Update/req
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1271_inst_ack_0, ack => ct_core_CP_34_elements(429)); -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(429), ack => WPIPE_ConvTranspose_output_pipe_1271_inst_req_1); -- 
    -- CP-element group 430:  transition  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	431 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_update_completed_
      -- CP-element group 430: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_Update/$exit
      -- CP-element group 430: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1271_Update/ack
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1271_inst_ack_1, ack => ct_core_CP_34_elements(430)); -- 
    -- CP-element group 431:  join  transition  output  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	411 
    -- CP-element group 431: 	430 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	432 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_sample_start_
      -- CP-element group 431: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_Sample/$entry
      -- CP-element group 431: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_Sample/req
      -- 
    req_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(431), ack => WPIPE_ConvTranspose_output_pipe_1274_inst_req_0); -- 
    ct_core_cp_element_group_431: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_431"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(411) & ct_core_CP_34_elements(430);
      gj_ct_core_cp_element_group_431 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(431), clk => clk, reset => reset); --
    end block;
    -- CP-element group 432:  transition  input  output  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	431 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	433 
    -- CP-element group 432:  members (6) 
      -- CP-element group 432: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_sample_completed_
      -- CP-element group 432: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_update_start_
      -- CP-element group 432: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_Sample/ack
      -- CP-element group 432: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_Update/$entry
      -- CP-element group 432: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_Update/req
      -- 
    ack_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1274_inst_ack_0, ack => ct_core_CP_34_elements(432)); -- 
    req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(432), ack => WPIPE_ConvTranspose_output_pipe_1274_inst_req_1); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	432 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	434 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_update_completed_
      -- CP-element group 433: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_Update/$exit
      -- CP-element group 433: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1274_Update/ack
      -- 
    ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1274_inst_ack_1, ack => ct_core_CP_34_elements(433)); -- 
    -- CP-element group 434:  join  transition  output  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	409 
    -- CP-element group 434: 	433 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	435 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_sample_start_
      -- CP-element group 434: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_Sample/$entry
      -- CP-element group 434: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_Sample/req
      -- 
    req_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(434), ack => WPIPE_ConvTranspose_output_pipe_1277_inst_req_0); -- 
    ct_core_cp_element_group_434: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_434"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(409) & ct_core_CP_34_elements(433);
      gj_ct_core_cp_element_group_434 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(434), clk => clk, reset => reset); --
    end block;
    -- CP-element group 435:  transition  input  output  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	434 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435:  members (6) 
      -- CP-element group 435: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_sample_completed_
      -- CP-element group 435: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_update_start_
      -- CP-element group 435: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_Sample/$exit
      -- CP-element group 435: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_Sample/ack
      -- CP-element group 435: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_Update/$entry
      -- CP-element group 435: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_Update/req
      -- 
    ack_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1277_inst_ack_0, ack => ct_core_CP_34_elements(435)); -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(435), ack => WPIPE_ConvTranspose_output_pipe_1277_inst_req_1); -- 
    -- CP-element group 436:  transition  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	435 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	437 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_update_completed_
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_Update/$exit
      -- CP-element group 436: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1277_Update/ack
      -- 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1277_inst_ack_1, ack => ct_core_CP_34_elements(436)); -- 
    -- CP-element group 437:  join  transition  output  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	407 
    -- CP-element group 437: 	436 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	438 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_sample_start_
      -- CP-element group 437: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_Sample/$entry
      -- CP-element group 437: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_Sample/req
      -- 
    req_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(437), ack => WPIPE_ConvTranspose_output_pipe_1280_inst_req_0); -- 
    ct_core_cp_element_group_437: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_437"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(407) & ct_core_CP_34_elements(436);
      gj_ct_core_cp_element_group_437 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(437), clk => clk, reset => reset); --
    end block;
    -- CP-element group 438:  transition  input  output  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	437 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	439 
    -- CP-element group 438:  members (6) 
      -- CP-element group 438: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_sample_completed_
      -- CP-element group 438: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_update_start_
      -- CP-element group 438: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_Sample/$exit
      -- CP-element group 438: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_Sample/ack
      -- CP-element group 438: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_Update/req
      -- 
    ack_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1280_inst_ack_0, ack => ct_core_CP_34_elements(438)); -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(438), ack => WPIPE_ConvTranspose_output_pipe_1280_inst_req_1); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	438 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	440 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_update_completed_
      -- CP-element group 439: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_Update/$exit
      -- CP-element group 439: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1280_Update/ack
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1280_inst_ack_1, ack => ct_core_CP_34_elements(439)); -- 
    -- CP-element group 440:  join  transition  output  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	405 
    -- CP-element group 440: 	439 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	441 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_sample_start_
      -- CP-element group 440: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_Sample/$entry
      -- CP-element group 440: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_Sample/req
      -- 
    req_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(440), ack => WPIPE_ConvTranspose_output_pipe_1283_inst_req_0); -- 
    ct_core_cp_element_group_440: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_440"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(405) & ct_core_CP_34_elements(439);
      gj_ct_core_cp_element_group_440 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(440), clk => clk, reset => reset); --
    end block;
    -- CP-element group 441:  transition  input  output  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	440 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	442 
    -- CP-element group 441:  members (6) 
      -- CP-element group 441: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_sample_completed_
      -- CP-element group 441: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_update_start_
      -- CP-element group 441: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_Sample/$exit
      -- CP-element group 441: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_Sample/ack
      -- CP-element group 441: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_Update/$entry
      -- CP-element group 441: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_Update/req
      -- 
    ack_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1283_inst_ack_0, ack => ct_core_CP_34_elements(441)); -- 
    req_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(441), ack => WPIPE_ConvTranspose_output_pipe_1283_inst_req_1); -- 
    -- CP-element group 442:  branch  transition  place  input  output  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	441 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	443 
    -- CP-element group 442: 	444 
    -- CP-element group 442:  members (17) 
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285__exit__
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_1292__entry__
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_1292__exit__
      -- CP-element group 442: 	 branch_block_stmt_25/if_stmt_1293__entry__
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/$exit
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_update_completed_
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_Update/$exit
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_1191_to_assign_stmt_1285/WPIPE_ConvTranspose_output_pipe_1283_Update/ack
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_1292/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/assign_stmt_1292/$exit
      -- CP-element group 442: 	 branch_block_stmt_25/if_stmt_1293_dead_link/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/if_stmt_1293_eval_test/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/if_stmt_1293_eval_test/$exit
      -- CP-element group 442: 	 branch_block_stmt_25/if_stmt_1293_eval_test/branch_req
      -- CP-element group 442: 	 branch_block_stmt_25/R_cmp264449_1294_place
      -- CP-element group 442: 	 branch_block_stmt_25/if_stmt_1293_if_link/$entry
      -- CP-element group 442: 	 branch_block_stmt_25/if_stmt_1293_else_link/$entry
      -- 
    ack_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1283_inst_ack_1, ack => ct_core_CP_34_elements(442)); -- 
    branch_req_2679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(442), ack => if_stmt_1293_branch_req_0); -- 
    -- CP-element group 443:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	442 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	445 
    -- CP-element group 443: 	446 
    -- CP-element group 443:  members (18) 
      -- CP-element group 443: 	 branch_block_stmt_25/merge_stmt_1299__exit__
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334__entry__
      -- CP-element group 443: 	 branch_block_stmt_25/if_stmt_1293_if_link/$exit
      -- CP-element group 443: 	 branch_block_stmt_25/if_stmt_1293_if_link/if_choice_transition
      -- CP-element group 443: 	 branch_block_stmt_25/forx_xend273_bbx_xnph
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_sample_start_
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_update_start_
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_Sample/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_Sample/rr
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_Update/cr
      -- CP-element group 443: 	 branch_block_stmt_25/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 443: 	 branch_block_stmt_25/merge_stmt_1299_PhiReqMerge
      -- CP-element group 443: 	 branch_block_stmt_25/merge_stmt_1299_PhiAck/$entry
      -- CP-element group 443: 	 branch_block_stmt_25/merge_stmt_1299_PhiAck/$exit
      -- CP-element group 443: 	 branch_block_stmt_25/merge_stmt_1299_PhiAck/dummy
      -- 
    if_choice_transition_2684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1293_branch_ack_1, ack => ct_core_CP_34_elements(443)); -- 
    rr_2701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(443), ack => type_cast_1320_inst_req_0); -- 
    cr_2706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(443), ack => type_cast_1320_inst_req_1); -- 
    -- CP-element group 444:  transition  place  input  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	442 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	522 
    -- CP-element group 444:  members (5) 
      -- CP-element group 444: 	 branch_block_stmt_25/if_stmt_1293_else_link/$exit
      -- CP-element group 444: 	 branch_block_stmt_25/if_stmt_1293_else_link/else_choice_transition
      -- CP-element group 444: 	 branch_block_stmt_25/forx_xend273_forx_xend444
      -- CP-element group 444: 	 branch_block_stmt_25/forx_xend273_forx_xend444_PhiReq/$entry
      -- CP-element group 444: 	 branch_block_stmt_25/forx_xend273_forx_xend444_PhiReq/$exit
      -- 
    else_choice_transition_2688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1293_branch_ack_0, ack => ct_core_CP_34_elements(444)); -- 
    -- CP-element group 445:  transition  input  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	443 
    -- CP-element group 445: successors 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_sample_completed_
      -- CP-element group 445: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_Sample/$exit
      -- CP-element group 445: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_Sample/ra
      -- 
    ra_2702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_0, ack => ct_core_CP_34_elements(445)); -- 
    -- CP-element group 446:  transition  place  input  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	443 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	516 
    -- CP-element group 446:  members (9) 
      -- CP-element group 446: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334__exit__
      -- CP-element group 446: 	 branch_block_stmt_25/bbx_xnph_forx_xbody371
      -- CP-element group 446: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/$exit
      -- CP-element group 446: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_update_completed_
      -- CP-element group 446: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_Update/$exit
      -- CP-element group 446: 	 branch_block_stmt_25/assign_stmt_1305_to_assign_stmt_1334/type_cast_1320_Update/ca
      -- CP-element group 446: 	 branch_block_stmt_25/bbx_xnph_forx_xbody371_PhiReq/$entry
      -- CP-element group 446: 	 branch_block_stmt_25/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1337/$entry
      -- CP-element group 446: 	 branch_block_stmt_25/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/$entry
      -- 
    ca_2707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1320_inst_ack_1, ack => ct_core_CP_34_elements(446)); -- 
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	521 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	492 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_final_index_sum_regn_sample_complete
      -- CP-element group 447: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_final_index_sum_regn_Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_final_index_sum_regn_Sample/ack
      -- 
    ack_2736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1349_index_offset_ack_0, ack => ct_core_CP_34_elements(447)); -- 
    -- CP-element group 448:  transition  input  output  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	521 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (11) 
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_sample_start_
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_root_address_calculated
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_offset_calculated
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_final_index_sum_regn_Update/$exit
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_final_index_sum_regn_Update/ack
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_base_plus_offset/$entry
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_base_plus_offset/$exit
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_base_plus_offset/sum_rename_req
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_base_plus_offset/sum_rename_ack
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_request/$entry
      -- CP-element group 448: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_request/req
      -- 
    ack_2741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1349_index_offset_ack_1, ack => ct_core_CP_34_elements(448)); -- 
    req_2750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(448), ack => addr_of_1350_final_reg_req_0); -- 
    -- CP-element group 449:  transition  input  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_sample_completed_
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_request/$exit
      -- CP-element group 449: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_request/ack
      -- 
    ack_2751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1350_final_reg_ack_0, ack => ct_core_CP_34_elements(449)); -- 
    -- CP-element group 450:  join  fork  transition  input  output  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	521 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (24) 
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_update_completed_
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_complete/$exit
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_complete/ack
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_sample_start_
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_base_address_calculated
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_word_address_calculated
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_root_address_calculated
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_base_address_resized
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_base_addr_resize/$entry
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_base_addr_resize/$exit
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_base_addr_resize/base_resize_req
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_base_addr_resize/base_resize_ack
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_base_plus_offset/$entry
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_base_plus_offset/$exit
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_base_plus_offset/sum_rename_req
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_base_plus_offset/sum_rename_ack
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_word_addrgen/$entry
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_word_addrgen/$exit
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_word_addrgen/root_register_req
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_word_addrgen/root_register_ack
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Sample/$entry
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Sample/word_access_start/$entry
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Sample/word_access_start/word_0/$entry
      -- CP-element group 450: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Sample/word_access_start/word_0/rr
      -- 
    ack_2756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1350_final_reg_ack_1, ack => ct_core_CP_34_elements(450)); -- 
    rr_2789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(450), ack => ptr_deref_1354_load_0_req_0); -- 
    -- CP-element group 451:  transition  input  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451:  members (5) 
      -- CP-element group 451: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_sample_completed_
      -- CP-element group 451: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Sample/$exit
      -- CP-element group 451: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Sample/word_access_start/$exit
      -- CP-element group 451: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Sample/word_access_start/word_0/$exit
      -- CP-element group 451: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Sample/word_access_start/word_0/ra
      -- 
    ra_2790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1354_load_0_ack_0, ack => ct_core_CP_34_elements(451)); -- 
    -- CP-element group 452:  fork  transition  input  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	521 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452: 	455 
    -- CP-element group 452: 	457 
    -- CP-element group 452: 	459 
    -- CP-element group 452: 	461 
    -- CP-element group 452: 	463 
    -- CP-element group 452: 	465 
    -- CP-element group 452: 	467 
    -- CP-element group 452:  members (33) 
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_update_completed_
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/$exit
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/word_access_complete/$exit
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/word_access_complete/word_0/$exit
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/word_access_complete/word_0/ca
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/ptr_deref_1354_Merge/$entry
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/ptr_deref_1354_Merge/$exit
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/ptr_deref_1354_Merge/merge_req
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/ptr_deref_1354_Merge/merge_ack
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_sample_start_
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_Sample/$entry
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_Sample/rr
      -- CP-element group 452: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_sample_start_
      -- 
    ca_2801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1354_load_0_ack_1, ack => ct_core_CP_34_elements(452)); -- 
    rr_2814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(452), ack => type_cast_1358_inst_req_0); -- 
    rr_2828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(452), ack => type_cast_1368_inst_req_0); -- 
    rr_2842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(452), ack => type_cast_1378_inst_req_0); -- 
    rr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(452), ack => type_cast_1388_inst_req_0); -- 
    rr_2870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(452), ack => type_cast_1398_inst_req_0); -- 
    rr_2884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(452), ack => type_cast_1408_inst_req_0); -- 
    rr_2898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(452), ack => type_cast_1418_inst_req_0); -- 
    rr_2912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(452), ack => type_cast_1428_inst_req_0); -- 
    -- CP-element group 453:  transition  input  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_sample_completed_
      -- CP-element group 453: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_Sample/$exit
      -- CP-element group 453: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_Sample/ra
      -- 
    ra_2815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_0, ack => ct_core_CP_34_elements(453)); -- 
    -- CP-element group 454:  transition  input  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	521 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	489 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_update_completed_
      -- CP-element group 454: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_Update/$exit
      -- CP-element group 454: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_Update/ca
      -- 
    ca_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_1, ack => ct_core_CP_34_elements(454)); -- 
    -- CP-element group 455:  transition  input  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	452 
    -- CP-element group 455: successors 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_Sample/ra
      -- CP-element group 455: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_Sample/$exit
      -- CP-element group 455: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_sample_completed_
      -- 
    ra_2829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_0, ack => ct_core_CP_34_elements(455)); -- 
    -- CP-element group 456:  transition  input  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	521 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	486 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_Update/$exit
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_Update/ca
      -- CP-element group 456: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_update_completed_
      -- 
    ca_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_1, ack => ct_core_CP_34_elements(456)); -- 
    -- CP-element group 457:  transition  input  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	452 
    -- CP-element group 457: successors 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_Sample/ra
      -- CP-element group 457: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_sample_completed_
      -- CP-element group 457: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_Sample/$exit
      -- 
    ra_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_0, ack => ct_core_CP_34_elements(457)); -- 
    -- CP-element group 458:  transition  input  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	521 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	483 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_Update/ca
      -- CP-element group 458: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_update_completed_
      -- CP-element group 458: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_Update/$exit
      -- 
    ca_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_1, ack => ct_core_CP_34_elements(458)); -- 
    -- CP-element group 459:  transition  input  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	452 
    -- CP-element group 459: successors 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_sample_completed_
      -- CP-element group 459: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_Sample/ra
      -- CP-element group 459: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_Sample/$exit
      -- 
    ra_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_0, ack => ct_core_CP_34_elements(459)); -- 
    -- CP-element group 460:  transition  input  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	521 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	480 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_Update/$exit
      -- CP-element group 460: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_Update/ca
      -- CP-element group 460: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_update_completed_
      -- 
    ca_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_1, ack => ct_core_CP_34_elements(460)); -- 
    -- CP-element group 461:  transition  input  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	452 
    -- CP-element group 461: successors 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_sample_completed_
      -- CP-element group 461: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_Sample/ra
      -- CP-element group 461: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_Sample/$exit
      -- 
    ra_2871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1398_inst_ack_0, ack => ct_core_CP_34_elements(461)); -- 
    -- CP-element group 462:  transition  input  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	521 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	477 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_Update/ca
      -- CP-element group 462: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_Update/$exit
      -- CP-element group 462: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_update_completed_
      -- 
    ca_2876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1398_inst_ack_1, ack => ct_core_CP_34_elements(462)); -- 
    -- CP-element group 463:  transition  input  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	452 
    -- CP-element group 463: successors 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_Sample/ra
      -- CP-element group 463: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_Sample/$exit
      -- CP-element group 463: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_sample_completed_
      -- 
    ra_2885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1408_inst_ack_0, ack => ct_core_CP_34_elements(463)); -- 
    -- CP-element group 464:  transition  input  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	521 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	474 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_Update/ca
      -- CP-element group 464: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_Update/$exit
      -- CP-element group 464: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_update_completed_
      -- 
    ca_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1408_inst_ack_1, ack => ct_core_CP_34_elements(464)); -- 
    -- CP-element group 465:  transition  input  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	452 
    -- CP-element group 465: successors 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_Sample/$exit
      -- CP-element group 465: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_Sample/ra
      -- CP-element group 465: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_sample_completed_
      -- 
    ra_2899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_0, ack => ct_core_CP_34_elements(465)); -- 
    -- CP-element group 466:  transition  input  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	521 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	471 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_Update/ca
      -- CP-element group 466: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_update_completed_
      -- CP-element group 466: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_Update/$exit
      -- 
    ca_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_1, ack => ct_core_CP_34_elements(466)); -- 
    -- CP-element group 467:  transition  input  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	452 
    -- CP-element group 467: successors 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_Sample/ra
      -- CP-element group 467: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_Sample/$exit
      -- CP-element group 467: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_sample_completed_
      -- 
    ra_2913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1428_inst_ack_0, ack => ct_core_CP_34_elements(467)); -- 
    -- CP-element group 468:  transition  input  output  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	521 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	469 
    -- CP-element group 468:  members (6) 
      -- CP-element group 468: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_update_completed_
      -- CP-element group 468: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_Sample/req
      -- CP-element group 468: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_Update/$exit
      -- CP-element group 468: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_Update/ca
      -- CP-element group 468: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_sample_start_
      -- CP-element group 468: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_Sample/$entry
      -- 
    ca_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1428_inst_ack_1, ack => ct_core_CP_34_elements(468)); -- 
    req_2926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(468), ack => WPIPE_ConvTranspose_output_pipe_1430_inst_req_0); -- 
    -- CP-element group 469:  transition  input  output  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	468 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	470 
    -- CP-element group 469:  members (6) 
      -- CP-element group 469: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_Sample/ack
      -- CP-element group 469: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_Sample/$exit
      -- CP-element group 469: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_Update/req
      -- CP-element group 469: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_Update/$entry
      -- CP-element group 469: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_sample_completed_
      -- CP-element group 469: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_update_start_
      -- 
    ack_2927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1430_inst_ack_0, ack => ct_core_CP_34_elements(469)); -- 
    req_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(469), ack => WPIPE_ConvTranspose_output_pipe_1430_inst_req_1); -- 
    -- CP-element group 470:  transition  input  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	469 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	471 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_Update/$exit
      -- CP-element group 470: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_Update/ack
      -- CP-element group 470: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1430_update_completed_
      -- 
    ack_2932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1430_inst_ack_1, ack => ct_core_CP_34_elements(470)); -- 
    -- CP-element group 471:  join  transition  output  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	466 
    -- CP-element group 471: 	470 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	472 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_sample_start_
      -- CP-element group 471: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_Sample/req
      -- CP-element group 471: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_Sample/$entry
      -- 
    req_2940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(471), ack => WPIPE_ConvTranspose_output_pipe_1433_inst_req_0); -- 
    ct_core_cp_element_group_471: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_471"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(466) & ct_core_CP_34_elements(470);
      gj_ct_core_cp_element_group_471 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(471), clk => clk, reset => reset); --
    end block;
    -- CP-element group 472:  transition  input  output  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	471 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	473 
    -- CP-element group 472:  members (6) 
      -- CP-element group 472: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_Update/req
      -- CP-element group 472: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_Update/$entry
      -- CP-element group 472: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_Sample/ack
      -- CP-element group 472: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_Sample/$exit
      -- CP-element group 472: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_update_start_
      -- CP-element group 472: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_sample_completed_
      -- 
    ack_2941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1433_inst_ack_0, ack => ct_core_CP_34_elements(472)); -- 
    req_2945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(472), ack => WPIPE_ConvTranspose_output_pipe_1433_inst_req_1); -- 
    -- CP-element group 473:  transition  input  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	472 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473:  members (3) 
      -- CP-element group 473: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_Update/ack
      -- CP-element group 473: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_Update/$exit
      -- CP-element group 473: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1433_update_completed_
      -- 
    ack_2946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1433_inst_ack_1, ack => ct_core_CP_34_elements(473)); -- 
    -- CP-element group 474:  join  transition  output  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	464 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474:  members (3) 
      -- CP-element group 474: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_Sample/req
      -- CP-element group 474: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_Sample/$entry
      -- CP-element group 474: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_sample_start_
      -- 
    req_2954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(474), ack => WPIPE_ConvTranspose_output_pipe_1436_inst_req_0); -- 
    ct_core_cp_element_group_474: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_474"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(464) & ct_core_CP_34_elements(473);
      gj_ct_core_cp_element_group_474 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(474), clk => clk, reset => reset); --
    end block;
    -- CP-element group 475:  transition  input  output  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	474 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	476 
    -- CP-element group 475:  members (6) 
      -- CP-element group 475: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_Update/req
      -- CP-element group 475: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_Sample/ack
      -- CP-element group 475: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_Sample/$exit
      -- CP-element group 475: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_update_start_
      -- CP-element group 475: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_sample_completed_
      -- 
    ack_2955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1436_inst_ack_0, ack => ct_core_CP_34_elements(475)); -- 
    req_2959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(475), ack => WPIPE_ConvTranspose_output_pipe_1436_inst_req_1); -- 
    -- CP-element group 476:  transition  input  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	475 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	477 
    -- CP-element group 476:  members (3) 
      -- CP-element group 476: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_Update/ack
      -- CP-element group 476: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_Update/$exit
      -- CP-element group 476: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1436_update_completed_
      -- 
    ack_2960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1436_inst_ack_1, ack => ct_core_CP_34_elements(476)); -- 
    -- CP-element group 477:  join  transition  output  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	462 
    -- CP-element group 477: 	476 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	478 
    -- CP-element group 477:  members (3) 
      -- CP-element group 477: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_Sample/req
      -- CP-element group 477: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_Sample/$entry
      -- CP-element group 477: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_sample_start_
      -- 
    req_2968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(477), ack => WPIPE_ConvTranspose_output_pipe_1439_inst_req_0); -- 
    ct_core_cp_element_group_477: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_477"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(462) & ct_core_CP_34_elements(476);
      gj_ct_core_cp_element_group_477 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(477), clk => clk, reset => reset); --
    end block;
    -- CP-element group 478:  transition  input  output  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	477 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	479 
    -- CP-element group 478:  members (6) 
      -- CP-element group 478: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_Update/req
      -- CP-element group 478: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_Sample/ack
      -- CP-element group 478: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_Sample/$exit
      -- CP-element group 478: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_update_start_
      -- CP-element group 478: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_sample_completed_
      -- 
    ack_2969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1439_inst_ack_0, ack => ct_core_CP_34_elements(478)); -- 
    req_2973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(478), ack => WPIPE_ConvTranspose_output_pipe_1439_inst_req_1); -- 
    -- CP-element group 479:  transition  input  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	478 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	480 
    -- CP-element group 479:  members (3) 
      -- CP-element group 479: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_Update/ack
      -- CP-element group 479: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_Update/$exit
      -- CP-element group 479: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1439_update_completed_
      -- 
    ack_2974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1439_inst_ack_1, ack => ct_core_CP_34_elements(479)); -- 
    -- CP-element group 480:  join  transition  output  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	460 
    -- CP-element group 480: 	479 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	481 
    -- CP-element group 480:  members (3) 
      -- CP-element group 480: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_Sample/req
      -- CP-element group 480: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_sample_start_
      -- CP-element group 480: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_Sample/$entry
      -- 
    req_2982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(480), ack => WPIPE_ConvTranspose_output_pipe_1442_inst_req_0); -- 
    ct_core_cp_element_group_480: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_480"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(460) & ct_core_CP_34_elements(479);
      gj_ct_core_cp_element_group_480 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(480), clk => clk, reset => reset); --
    end block;
    -- CP-element group 481:  transition  input  output  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	480 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	482 
    -- CP-element group 481:  members (6) 
      -- CP-element group 481: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_sample_completed_
      -- CP-element group 481: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_Update/req
      -- CP-element group 481: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_update_start_
      -- CP-element group 481: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_Sample/ack
      -- CP-element group 481: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_Sample/$exit
      -- 
    ack_2983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1442_inst_ack_0, ack => ct_core_CP_34_elements(481)); -- 
    req_2987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(481), ack => WPIPE_ConvTranspose_output_pipe_1442_inst_req_1); -- 
    -- CP-element group 482:  transition  input  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	481 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	483 
    -- CP-element group 482:  members (3) 
      -- CP-element group 482: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_Update/$exit
      -- CP-element group 482: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_update_completed_
      -- CP-element group 482: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1442_Update/ack
      -- 
    ack_2988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1442_inst_ack_1, ack => ct_core_CP_34_elements(482)); -- 
    -- CP-element group 483:  join  transition  output  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	458 
    -- CP-element group 483: 	482 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	484 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_Sample/req
      -- CP-element group 483: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_Sample/$entry
      -- CP-element group 483: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_sample_start_
      -- 
    req_2996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(483), ack => WPIPE_ConvTranspose_output_pipe_1445_inst_req_0); -- 
    ct_core_cp_element_group_483: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_483"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(458) & ct_core_CP_34_elements(482);
      gj_ct_core_cp_element_group_483 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(483), clk => clk, reset => reset); --
    end block;
    -- CP-element group 484:  transition  input  output  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	483 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	485 
    -- CP-element group 484:  members (6) 
      -- CP-element group 484: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_Update/$entry
      -- CP-element group 484: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_Update/req
      -- CP-element group 484: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_Sample/$exit
      -- CP-element group 484: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_Sample/ack
      -- CP-element group 484: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_sample_completed_
      -- CP-element group 484: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_update_start_
      -- 
    ack_2997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1445_inst_ack_0, ack => ct_core_CP_34_elements(484)); -- 
    req_3001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(484), ack => WPIPE_ConvTranspose_output_pipe_1445_inst_req_1); -- 
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	484 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	486 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_Update/$exit
      -- CP-element group 485: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_Update/ack
      -- CP-element group 485: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1445_update_completed_
      -- 
    ack_3002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1445_inst_ack_1, ack => ct_core_CP_34_elements(485)); -- 
    -- CP-element group 486:  join  transition  output  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	456 
    -- CP-element group 486: 	485 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (3) 
      -- CP-element group 486: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_sample_start_
      -- CP-element group 486: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_Sample/$entry
      -- CP-element group 486: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_Sample/req
      -- 
    req_3010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(486), ack => WPIPE_ConvTranspose_output_pipe_1448_inst_req_0); -- 
    ct_core_cp_element_group_486: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_486"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(456) & ct_core_CP_34_elements(485);
      gj_ct_core_cp_element_group_486 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(486), clk => clk, reset => reset); --
    end block;
    -- CP-element group 487:  transition  input  output  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	488 
    -- CP-element group 487:  members (6) 
      -- CP-element group 487: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_sample_completed_
      -- CP-element group 487: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_update_start_
      -- CP-element group 487: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_Sample/$exit
      -- CP-element group 487: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_Sample/ack
      -- CP-element group 487: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_Update/$entry
      -- CP-element group 487: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_Update/req
      -- 
    ack_3011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0, ack => ct_core_CP_34_elements(487)); -- 
    req_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(487), ack => WPIPE_ConvTranspose_output_pipe_1448_inst_req_1); -- 
    -- CP-element group 488:  transition  input  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	487 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	489 
    -- CP-element group 488:  members (3) 
      -- CP-element group 488: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_update_completed_
      -- CP-element group 488: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_Update/ack
      -- CP-element group 488: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1448_Update/$exit
      -- 
    ack_3016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1, ack => ct_core_CP_34_elements(488)); -- 
    -- CP-element group 489:  join  transition  output  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	454 
    -- CP-element group 489: 	488 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	490 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_Sample/req
      -- CP-element group 489: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_sample_start_
      -- 
    req_3024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(489), ack => WPIPE_ConvTranspose_output_pipe_1451_inst_req_0); -- 
    ct_core_cp_element_group_489: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_489"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(454) & ct_core_CP_34_elements(488);
      gj_ct_core_cp_element_group_489 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(489), clk => clk, reset => reset); --
    end block;
    -- CP-element group 490:  transition  input  output  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	489 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	491 
    -- CP-element group 490:  members (6) 
      -- CP-element group 490: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_Sample/ack
      -- CP-element group 490: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_Sample/$exit
      -- CP-element group 490: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_Update/$entry
      -- CP-element group 490: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_Update/req
      -- CP-element group 490: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_update_start_
      -- CP-element group 490: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_sample_completed_
      -- 
    ack_3025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 490_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0, ack => ct_core_CP_34_elements(490)); -- 
    req_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(490), ack => WPIPE_ConvTranspose_output_pipe_1451_inst_req_1); -- 
    -- CP-element group 491:  transition  input  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	490 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	492 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_Update/$exit
      -- CP-element group 491: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_update_completed_
      -- CP-element group 491: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/WPIPE_ConvTranspose_output_pipe_1451_Update/ack
      -- 
    ack_3030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1, ack => ct_core_CP_34_elements(491)); -- 
    -- CP-element group 492:  branch  join  transition  place  output  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	447 
    -- CP-element group 492: 	491 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492: 	494 
    -- CP-element group 492:  members (10) 
      -- CP-element group 492: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464__exit__
      -- CP-element group 492: 	 branch_block_stmt_25/if_stmt_1465__entry__
      -- CP-element group 492: 	 branch_block_stmt_25/if_stmt_1465_dead_link/$entry
      -- CP-element group 492: 	 branch_block_stmt_25/if_stmt_1465_eval_test/$entry
      -- CP-element group 492: 	 branch_block_stmt_25/if_stmt_1465_eval_test/$exit
      -- CP-element group 492: 	 branch_block_stmt_25/if_stmt_1465_eval_test/branch_req
      -- CP-element group 492: 	 branch_block_stmt_25/if_stmt_1465_if_link/$entry
      -- CP-element group 492: 	 branch_block_stmt_25/R_exitcond1_1466_place
      -- CP-element group 492: 	 branch_block_stmt_25/if_stmt_1465_else_link/$entry
      -- CP-element group 492: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/$exit
      -- 
    branch_req_3038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(492), ack => if_stmt_1465_branch_req_0); -- 
    ct_core_cp_element_group_492: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_492"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(447) & ct_core_CP_34_elements(491);
      gj_ct_core_cp_element_group_492 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(492), clk => clk, reset => reset); --
    end block;
    -- CP-element group 493:  merge  transition  place  input  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	492 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	522 
    -- CP-element group 493:  members (13) 
      -- CP-element group 493: 	 branch_block_stmt_25/merge_stmt_1471__exit__
      -- CP-element group 493: 	 branch_block_stmt_25/forx_xend444x_xloopexit_forx_xend444
      -- CP-element group 493: 	 branch_block_stmt_25/if_stmt_1465_if_link/$exit
      -- CP-element group 493: 	 branch_block_stmt_25/if_stmt_1465_if_link/if_choice_transition
      -- CP-element group 493: 	 branch_block_stmt_25/forx_xbody371_forx_xend444x_xloopexit
      -- CP-element group 493: 	 branch_block_stmt_25/forx_xbody371_forx_xend444x_xloopexit_PhiReq/$entry
      -- CP-element group 493: 	 branch_block_stmt_25/forx_xbody371_forx_xend444x_xloopexit_PhiReq/$exit
      -- CP-element group 493: 	 branch_block_stmt_25/merge_stmt_1471_PhiReqMerge
      -- CP-element group 493: 	 branch_block_stmt_25/merge_stmt_1471_PhiAck/$entry
      -- CP-element group 493: 	 branch_block_stmt_25/merge_stmt_1471_PhiAck/$exit
      -- CP-element group 493: 	 branch_block_stmt_25/merge_stmt_1471_PhiAck/dummy
      -- CP-element group 493: 	 branch_block_stmt_25/forx_xend444x_xloopexit_forx_xend444_PhiReq/$entry
      -- CP-element group 493: 	 branch_block_stmt_25/forx_xend444x_xloopexit_forx_xend444_PhiReq/$exit
      -- 
    if_choice_transition_3043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1465_branch_ack_1, ack => ct_core_CP_34_elements(493)); -- 
    -- CP-element group 494:  fork  transition  place  input  output  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	492 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	517 
    -- CP-element group 494: 	518 
    -- CP-element group 494:  members (12) 
      -- CP-element group 494: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371
      -- CP-element group 494: 	 branch_block_stmt_25/if_stmt_1465_else_link/else_choice_transition
      -- CP-element group 494: 	 branch_block_stmt_25/if_stmt_1465_else_link/$exit
      -- CP-element group 494: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/$entry
      -- CP-element group 494: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/$entry
      -- CP-element group 494: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/$entry
      -- CP-element group 494: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/$entry
      -- CP-element group 494: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/SplitProtocol/$entry
      -- CP-element group 494: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/SplitProtocol/Sample/$entry
      -- CP-element group 494: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/SplitProtocol/Sample/rr
      -- CP-element group 494: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/SplitProtocol/Update/$entry
      -- CP-element group 494: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1465_branch_ack_0, ack => ct_core_CP_34_elements(494)); -- 
    rr_3322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(494), ack => type_cast_1343_inst_req_0); -- 
    cr_3327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(494), ack => type_cast_1343_inst_req_1); -- 
    -- CP-element group 495:  merge  branch  transition  place  output  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	118 
    -- CP-element group 495: 	163 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	119 
    -- CP-element group 495: 	120 
    -- CP-element group 495:  members (17) 
      -- CP-element group 495: 	 branch_block_stmt_25/merge_stmt_401__exit__
      -- CP-element group 495: 	 branch_block_stmt_25/assign_stmt_407__entry__
      -- CP-element group 495: 	 branch_block_stmt_25/assign_stmt_407__exit__
      -- CP-element group 495: 	 branch_block_stmt_25/if_stmt_408__entry__
      -- CP-element group 495: 	 branch_block_stmt_25/assign_stmt_407/$entry
      -- CP-element group 495: 	 branch_block_stmt_25/assign_stmt_407/$exit
      -- CP-element group 495: 	 branch_block_stmt_25/if_stmt_408_dead_link/$entry
      -- CP-element group 495: 	 branch_block_stmt_25/if_stmt_408_eval_test/$entry
      -- CP-element group 495: 	 branch_block_stmt_25/if_stmt_408_eval_test/$exit
      -- CP-element group 495: 	 branch_block_stmt_25/if_stmt_408_eval_test/branch_req
      -- CP-element group 495: 	 branch_block_stmt_25/R_cmp175463_409_place
      -- CP-element group 495: 	 branch_block_stmt_25/if_stmt_408_if_link/$entry
      -- CP-element group 495: 	 branch_block_stmt_25/if_stmt_408_else_link/$entry
      -- CP-element group 495: 	 branch_block_stmt_25/merge_stmt_401_PhiAck/dummy
      -- CP-element group 495: 	 branch_block_stmt_25/merge_stmt_401_PhiAck/$exit
      -- CP-element group 495: 	 branch_block_stmt_25/merge_stmt_401_PhiAck/$entry
      -- CP-element group 495: 	 branch_block_stmt_25/merge_stmt_401_PhiReqMerge
      -- 
    branch_req_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(495), ack => if_stmt_408_branch_req_0); -- 
    ct_core_CP_34_elements(495) <= OrReduce(ct_core_CP_34_elements(118) & ct_core_CP_34_elements(163));
    -- CP-element group 496:  transition  output  delay-element  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	122 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	500 
    -- CP-element group 496:  members (5) 
      -- CP-element group 496: 	 branch_block_stmt_25/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_req
      -- CP-element group 496: 	 branch_block_stmt_25/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_456_konst_delay_trans
      -- CP-element group 496: 	 branch_block_stmt_25/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/$exit
      -- CP-element group 496: 	 branch_block_stmt_25/bbx_xnph469_forx_xbody_PhiReq/phi_stmt_452/$exit
      -- CP-element group 496: 	 branch_block_stmt_25/bbx_xnph469_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_452_req_3095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_452_req_3095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(496), ack => phi_stmt_452_req_0); -- 
    -- Element group ct_core_CP_34_elements(496) is a control-delay.
    cp_element_496_delay: control_delay_element  generic map(name => " 496_delay", delay_value => 1)  port map(req => ct_core_CP_34_elements(122), ack => ct_core_CP_34_elements(496), clk => clk, reset =>reset);
    -- CP-element group 497:  transition  input  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	164 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	499 
    -- CP-element group 497:  members (2) 
      -- CP-element group 497: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/SplitProtocol/Sample/$exit
      -- CP-element group 497: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/SplitProtocol/Sample/ra
      -- 
    ra_3115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 497_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_458_inst_ack_0, ack => ct_core_CP_34_elements(497)); -- 
    -- CP-element group 498:  transition  input  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	164 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	499 
    -- CP-element group 498:  members (2) 
      -- CP-element group 498: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/SplitProtocol/Update/ca
      -- CP-element group 498: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/SplitProtocol/Update/$exit
      -- 
    ca_3120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_458_inst_ack_1, ack => ct_core_CP_34_elements(498)); -- 
    -- CP-element group 499:  join  transition  output  bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	497 
    -- CP-element group 499: 	498 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	500 
    -- CP-element group 499:  members (6) 
      -- CP-element group 499: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/SplitProtocol/$exit
      -- CP-element group 499: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/$exit
      -- CP-element group 499: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/$exit
      -- CP-element group 499: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 499: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_sources/type_cast_458/$exit
      -- CP-element group 499: 	 branch_block_stmt_25/forx_xbody_forx_xbody_PhiReq/phi_stmt_452/phi_stmt_452_req
      -- 
    phi_stmt_452_req_3121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_452_req_3121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(499), ack => phi_stmt_452_req_1); -- 
    ct_core_cp_element_group_499: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_499"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(497) & ct_core_CP_34_elements(498);
      gj_ct_core_cp_element_group_499 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(499), clk => clk, reset => reset); --
    end block;
    -- CP-element group 500:  merge  transition  place  bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	496 
    -- CP-element group 500: 	499 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	501 
    -- CP-element group 500:  members (2) 
      -- CP-element group 500: 	 branch_block_stmt_25/merge_stmt_451_PhiReqMerge
      -- CP-element group 500: 	 branch_block_stmt_25/merge_stmt_451_PhiAck/$entry
      -- 
    ct_core_CP_34_elements(500) <= OrReduce(ct_core_CP_34_elements(496) & ct_core_CP_34_elements(499));
    -- CP-element group 501:  fork  transition  place  input  output  bypass 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	500 
    -- CP-element group 501: successors 
    -- CP-element group 501: 	123 
    -- CP-element group 501: 	124 
    -- CP-element group 501: 	126 
    -- CP-element group 501: 	127 
    -- CP-element group 501: 	130 
    -- CP-element group 501: 	134 
    -- CP-element group 501: 	138 
    -- CP-element group 501: 	142 
    -- CP-element group 501: 	146 
    -- CP-element group 501: 	150 
    -- CP-element group 501: 	154 
    -- CP-element group 501: 	158 
    -- CP-element group 501: 	161 
    -- CP-element group 501:  members (56) 
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_scale_1/scale_rename_req
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_scale_1/$exit
      -- CP-element group 501: 	 branch_block_stmt_25/merge_stmt_451__exit__
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614__entry__
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_update_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_final_index_sum_regn_Sample/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_final_index_sum_regn_Update/req
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_final_index_sum_regn_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_scale_1/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_final_index_sum_regn_Sample/req
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_resize_1/index_resize_ack
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_Update/cr
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_final_index_sum_regn_update_start
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_485_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_Update/cr
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Update/word_access_complete/word_0/cr
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Update/word_access_complete/word_0/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_scale_1/scale_rename_ack
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_resize_1/index_resize_req
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Update/word_access_complete/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_539_update_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_Update/cr
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_complete/req
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_Update/cr
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_Update/cr
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_Update/cr
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_Update/cr
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_472_update_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_557_update_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/ptr_deref_601_update_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_575_update_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_503_update_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_Update/cr
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_Sample/rr
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_Sample/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_521_update_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/RPIPE_ConvTranspose_input_pipe_468_sample_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_resize_1/$exit
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_resize_1/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_computed_1
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_complete/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/type_cast_593_update_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_scaled_1
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/$entry
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/addr_of_465_update_start_
      -- CP-element group 501: 	 branch_block_stmt_25/assign_stmt_466_to_assign_stmt_614/array_obj_ref_464_index_resized_1
      -- CP-element group 501: 	 branch_block_stmt_25/merge_stmt_451_PhiAck/phi_stmt_452_ack
      -- CP-element group 501: 	 branch_block_stmt_25/merge_stmt_451_PhiAck/$exit
      -- 
    phi_stmt_452_ack_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_452_ack_0, ack => ct_core_CP_34_elements(501)); -- 
    req_975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => array_obj_ref_464_index_offset_req_1); -- 
    req_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => array_obj_ref_464_index_offset_req_0); -- 
    cr_1046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => type_cast_485_inst_req_1); -- 
    cr_1130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => type_cast_539_inst_req_1); -- 
    cr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => ptr_deref_601_store_0_req_1); -- 
    cr_1074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => type_cast_503_inst_req_1); -- 
    req_990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => addr_of_465_final_reg_req_1); -- 
    cr_1214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => type_cast_593_inst_req_1); -- 
    cr_1018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => type_cast_472_inst_req_1); -- 
    cr_1158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => type_cast_557_inst_req_1); -- 
    cr_1186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => type_cast_575_inst_req_1); -- 
    cr_1102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => type_cast_521_inst_req_1); -- 
    rr_999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(501), ack => RPIPE_ConvTranspose_input_pipe_468_inst_req_0); -- 
    -- CP-element group 502:  transition  output  delay-element  bypass 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	166 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	506 
    -- CP-element group 502:  members (5) 
      -- CP-element group 502: 	 branch_block_stmt_25/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_req
      -- CP-element group 502: 	 branch_block_stmt_25/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_663_konst_delay_trans
      -- CP-element group 502: 	 branch_block_stmt_25/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/$exit
      -- CP-element group 502: 	 branch_block_stmt_25/bbx_xnph465_forx_xbody177_PhiReq/phi_stmt_659/$exit
      -- CP-element group 502: 	 branch_block_stmt_25/bbx_xnph465_forx_xbody177_PhiReq/$exit
      -- 
    phi_stmt_659_req_3149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_659_req_3149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(502), ack => phi_stmt_659_req_0); -- 
    -- Element group ct_core_CP_34_elements(502) is a control-delay.
    cp_element_502_delay: control_delay_element  generic map(name => " 502_delay", delay_value => 1)  port map(req => ct_core_CP_34_elements(166), ack => ct_core_CP_34_elements(502), clk => clk, reset =>reset);
    -- CP-element group 503:  transition  input  bypass 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	208 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	505 
    -- CP-element group 503:  members (2) 
      -- CP-element group 503: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/SplitProtocol/Sample/$exit
      -- CP-element group 503: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/SplitProtocol/Sample/ra
      -- 
    ra_3169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 503_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_665_inst_ack_0, ack => ct_core_CP_34_elements(503)); -- 
    -- CP-element group 504:  transition  input  bypass 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	208 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	505 
    -- CP-element group 504:  members (2) 
      -- CP-element group 504: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/SplitProtocol/Update/$exit
      -- CP-element group 504: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/SplitProtocol/Update/ca
      -- 
    ca_3174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_665_inst_ack_1, ack => ct_core_CP_34_elements(504)); -- 
    -- CP-element group 505:  join  transition  output  bypass 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	503 
    -- CP-element group 505: 	504 
    -- CP-element group 505: successors 
    -- CP-element group 505: 	506 
    -- CP-element group 505:  members (6) 
      -- CP-element group 505: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/$exit
      -- CP-element group 505: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/type_cast_665/SplitProtocol/$exit
      -- CP-element group 505: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_sources/$exit
      -- CP-element group 505: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/$exit
      -- CP-element group 505: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/phi_stmt_659/phi_stmt_659_req
      -- CP-element group 505: 	 branch_block_stmt_25/forx_xbody177_forx_xbody177_PhiReq/$exit
      -- 
    phi_stmt_659_req_3175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_659_req_3175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(505), ack => phi_stmt_659_req_1); -- 
    ct_core_cp_element_group_505: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_505"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(503) & ct_core_CP_34_elements(504);
      gj_ct_core_cp_element_group_505 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(505), clk => clk, reset => reset); --
    end block;
    -- CP-element group 506:  merge  transition  place  bypass 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	502 
    -- CP-element group 506: 	505 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	507 
    -- CP-element group 506:  members (2) 
      -- CP-element group 506: 	 branch_block_stmt_25/merge_stmt_658_PhiAck/$entry
      -- CP-element group 506: 	 branch_block_stmt_25/merge_stmt_658_PhiReqMerge
      -- 
    ct_core_CP_34_elements(506) <= OrReduce(ct_core_CP_34_elements(502) & ct_core_CP_34_elements(505));
    -- CP-element group 507:  fork  transition  place  input  output  bypass 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	506 
    -- CP-element group 507: successors 
    -- CP-element group 507: 	167 
    -- CP-element group 507: 	168 
    -- CP-element group 507: 	170 
    -- CP-element group 507: 	171 
    -- CP-element group 507: 	174 
    -- CP-element group 507: 	178 
    -- CP-element group 507: 	182 
    -- CP-element group 507: 	186 
    -- CP-element group 507: 	190 
    -- CP-element group 507: 	194 
    -- CP-element group 507: 	198 
    -- CP-element group 507: 	202 
    -- CP-element group 507: 	205 
    -- CP-element group 507:  members (56) 
      -- CP-element group 507: 	 branch_block_stmt_25/merge_stmt_658__exit__
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821__entry__
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_final_index_sum_regn_Update/req
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_Update/cr
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_final_index_sum_regn_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_complete/req
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_final_index_sum_regn_Sample/req
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_final_index_sum_regn_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_final_index_sum_regn_update_start
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_complete/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_scale_1/scale_rename_ack
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_Update/cr
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_scale_1/scale_rename_req
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_scale_1/$exit
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_scale_1/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_update_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_resize_1/index_resize_ack
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_resize_1/index_resize_req
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_679_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_resize_1/$exit
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_resize_1/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_Sample/rr
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_computed_1
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_scaled_1
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/array_obj_ref_671_index_resized_1
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/addr_of_672_update_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_692_update_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/RPIPE_ConvTranspose_input_pipe_675_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_update_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_710_Update/cr
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_update_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_728_Update/cr
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_update_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_746_Update/cr
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_update_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_764_Update/cr
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_update_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_782_Update/cr
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_update_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/type_cast_800_Update/cr
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_update_start_
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Update/word_access_complete/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Update/word_access_complete/word_0/$entry
      -- CP-element group 507: 	 branch_block_stmt_25/assign_stmt_673_to_assign_stmt_821/ptr_deref_808_Update/word_access_complete/word_0/cr
      -- CP-element group 507: 	 branch_block_stmt_25/merge_stmt_658_PhiAck/$exit
      -- CP-element group 507: 	 branch_block_stmt_25/merge_stmt_658_PhiAck/phi_stmt_659_ack
      -- 
    phi_stmt_659_ack_3180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 507_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_659_ack_0, ack => ct_core_CP_34_elements(507)); -- 
    req_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => array_obj_ref_671_index_offset_req_1); -- 
    cr_1405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => type_cast_692_inst_req_1); -- 
    req_1349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => addr_of_672_final_reg_req_1); -- 
    req_1329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => array_obj_ref_671_index_offset_req_0); -- 
    cr_1377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => type_cast_679_inst_req_1); -- 
    rr_1358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => RPIPE_ConvTranspose_input_pipe_675_inst_req_0); -- 
    cr_1433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => type_cast_710_inst_req_1); -- 
    cr_1461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => type_cast_728_inst_req_1); -- 
    cr_1489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => type_cast_746_inst_req_1); -- 
    cr_1517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => type_cast_764_inst_req_1); -- 
    cr_1545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => type_cast_782_inst_req_1); -- 
    cr_1573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => type_cast_800_inst_req_1); -- 
    cr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(507), ack => ptr_deref_808_store_0_req_1); -- 
    -- CP-element group 508:  merge  branch  transition  place  output  bypass 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	120 
    -- CP-element group 508: 	207 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	209 
    -- CP-element group 508: 	210 
    -- CP-element group 508:  members (17) 
      -- CP-element group 508: 	 branch_block_stmt_25/merge_stmt_830__exit__
      -- CP-element group 508: 	 branch_block_stmt_25/assign_stmt_836__entry__
      -- CP-element group 508: 	 branch_block_stmt_25/assign_stmt_836__exit__
      -- CP-element group 508: 	 branch_block_stmt_25/if_stmt_837__entry__
      -- CP-element group 508: 	 branch_block_stmt_25/merge_stmt_830_PhiReqMerge
      -- CP-element group 508: 	 branch_block_stmt_25/merge_stmt_830_PhiAck/$exit
      -- CP-element group 508: 	 branch_block_stmt_25/merge_stmt_830_PhiAck/dummy
      -- CP-element group 508: 	 branch_block_stmt_25/assign_stmt_836/$entry
      -- CP-element group 508: 	 branch_block_stmt_25/assign_stmt_836/$exit
      -- CP-element group 508: 	 branch_block_stmt_25/if_stmt_837_dead_link/$entry
      -- CP-element group 508: 	 branch_block_stmt_25/if_stmt_837_eval_test/$entry
      -- CP-element group 508: 	 branch_block_stmt_25/if_stmt_837_eval_test/$exit
      -- CP-element group 508: 	 branch_block_stmt_25/if_stmt_837_eval_test/branch_req
      -- CP-element group 508: 	 branch_block_stmt_25/R_cmp264448_838_place
      -- CP-element group 508: 	 branch_block_stmt_25/if_stmt_837_if_link/$entry
      -- CP-element group 508: 	 branch_block_stmt_25/if_stmt_837_else_link/$entry
      -- CP-element group 508: 	 branch_block_stmt_25/merge_stmt_830_PhiAck/$entry
      -- 
    branch_req_1654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(508), ack => if_stmt_837_branch_req_0); -- 
    ct_core_CP_34_elements(508) <= OrReduce(ct_core_CP_34_elements(120) & ct_core_CP_34_elements(207));
    -- CP-element group 509:  transition  output  delay-element  bypass 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	212 
    -- CP-element group 509: successors 
    -- CP-element group 509: 	513 
    -- CP-element group 509:  members (5) 
      -- CP-element group 509: 	 branch_block_stmt_25/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_req
      -- CP-element group 509: 	 branch_block_stmt_25/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/$exit
      -- CP-element group 509: 	 branch_block_stmt_25/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_885_konst_delay_trans
      -- CP-element group 509: 	 branch_block_stmt_25/bbx_xnph451_forx_xbody266_PhiReq/phi_stmt_881/$exit
      -- CP-element group 509: 	 branch_block_stmt_25/bbx_xnph451_forx_xbody266_PhiReq/$exit
      -- 
    phi_stmt_881_req_3226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_881_req_3226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(509), ack => phi_stmt_881_req_0); -- 
    -- Element group ct_core_CP_34_elements(509) is a control-delay.
    cp_element_509_delay: control_delay_element  generic map(name => " 509_delay", delay_value => 1)  port map(req => ct_core_CP_34_elements(212), ack => ct_core_CP_34_elements(509), clk => clk, reset =>reset);
    -- CP-element group 510:  transition  input  bypass 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	221 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	512 
    -- CP-element group 510:  members (2) 
      -- CP-element group 510: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/SplitProtocol/Sample/ra
      -- CP-element group 510: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/SplitProtocol/Sample/$exit
      -- 
    ra_3246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_0, ack => ct_core_CP_34_elements(510)); -- 
    -- CP-element group 511:  transition  input  bypass 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	221 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	512 
    -- CP-element group 511:  members (2) 
      -- CP-element group 511: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/SplitProtocol/Update/ca
      -- CP-element group 511: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/SplitProtocol/Update/$exit
      -- 
    ca_3251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 511_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_1, ack => ct_core_CP_34_elements(511)); -- 
    -- CP-element group 512:  join  transition  output  bypass 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	510 
    -- CP-element group 512: 	511 
    -- CP-element group 512: successors 
    -- CP-element group 512: 	513 
    -- CP-element group 512:  members (6) 
      -- CP-element group 512: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_req
      -- CP-element group 512: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/$exit
      -- CP-element group 512: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 512: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/SplitProtocol/$exit
      -- CP-element group 512: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/type_cast_887/$exit
      -- CP-element group 512: 	 branch_block_stmt_25/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_881/phi_stmt_881_sources/$exit
      -- 
    phi_stmt_881_req_3252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_881_req_3252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(512), ack => phi_stmt_881_req_1); -- 
    ct_core_cp_element_group_512: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_512"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(510) & ct_core_CP_34_elements(511);
      gj_ct_core_cp_element_group_512 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(512), clk => clk, reset => reset); --
    end block;
    -- CP-element group 513:  merge  transition  place  bypass 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	509 
    -- CP-element group 513: 	512 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	514 
    -- CP-element group 513:  members (2) 
      -- CP-element group 513: 	 branch_block_stmt_25/merge_stmt_880_PhiReqMerge
      -- CP-element group 513: 	 branch_block_stmt_25/merge_stmt_880_PhiAck/$entry
      -- 
    ct_core_CP_34_elements(513) <= OrReduce(ct_core_CP_34_elements(509) & ct_core_CP_34_elements(512));
    -- CP-element group 514:  fork  transition  place  input  output  bypass 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	513 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	218 
    -- CP-element group 514: 	213 
    -- CP-element group 514: 	214 
    -- CP-element group 514: 	216 
    -- CP-element group 514:  members (29) 
      -- CP-element group 514: 	 branch_block_stmt_25/merge_stmt_880__exit__
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911__entry__
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/$entry
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_update_start_
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_resized_1
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_scaled_1
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_computed_1
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_resize_1/$entry
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_resize_1/$exit
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_resize_1/index_resize_req
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_resize_1/index_resize_ack
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_scale_1/$entry
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_scale_1/$exit
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_scale_1/scale_rename_req
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_index_scale_1/scale_rename_ack
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_final_index_sum_regn_update_start
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_final_index_sum_regn_Sample/$entry
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_final_index_sum_regn_Sample/req
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_final_index_sum_regn_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/array_obj_ref_893_final_index_sum_regn_Update/req
      -- CP-element group 514: 	 branch_block_stmt_25/merge_stmt_880_PhiAck/phi_stmt_881_ack
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_complete/$entry
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/addr_of_894_complete/req
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_update_start_
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Update/word_access_complete/$entry
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Update/word_access_complete/word_0/$entry
      -- CP-element group 514: 	 branch_block_stmt_25/assign_stmt_895_to_assign_stmt_911/ptr_deref_897_Update/word_access_complete/word_0/cr
      -- CP-element group 514: 	 branch_block_stmt_25/merge_stmt_880_PhiAck/$exit
      -- 
    phi_stmt_881_ack_3257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_881_ack_0, ack => ct_core_CP_34_elements(514)); -- 
    req_1710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(514), ack => array_obj_ref_893_index_offset_req_0); -- 
    req_1715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(514), ack => array_obj_ref_893_index_offset_req_1); -- 
    req_1730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(514), ack => addr_of_894_final_reg_req_1); -- 
    cr_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(514), ack => ptr_deref_897_store_0_req_1); -- 
    -- CP-element group 515:  merge  fork  transition  place  output  bypass 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	220 
    -- CP-element group 515: 	210 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	222 
    -- CP-element group 515: 	223 
    -- CP-element group 515:  members (13) 
      -- CP-element group 515: 	 branch_block_stmt_25/merge_stmt_920__exit__
      -- CP-element group 515: 	 branch_block_stmt_25/call_stmt_923__entry__
      -- CP-element group 515: 	 branch_block_stmt_25/call_stmt_923/$entry
      -- CP-element group 515: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_sample_start_
      -- CP-element group 515: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_update_start_
      -- CP-element group 515: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_Sample/$entry
      -- CP-element group 515: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_Sample/crr
      -- CP-element group 515: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_Update/$entry
      -- CP-element group 515: 	 branch_block_stmt_25/call_stmt_923/call_stmt_923_Update/ccr
      -- CP-element group 515: 	 branch_block_stmt_25/merge_stmt_920_PhiReqMerge
      -- CP-element group 515: 	 branch_block_stmt_25/merge_stmt_920_PhiAck/$entry
      -- CP-element group 515: 	 branch_block_stmt_25/merge_stmt_920_PhiAck/$exit
      -- CP-element group 515: 	 branch_block_stmt_25/merge_stmt_920_PhiAck/dummy
      -- 
    crr_1811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(515), ack => call_stmt_923_call_req_0); -- 
    ccr_1816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(515), ack => call_stmt_923_call_req_1); -- 
    ct_core_CP_34_elements(515) <= OrReduce(ct_core_CP_34_elements(220) & ct_core_CP_34_elements(210));
    -- CP-element group 516:  transition  output  delay-element  bypass 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	446 
    -- CP-element group 516: successors 
    -- CP-element group 516: 	520 
    -- CP-element group 516:  members (5) 
      -- CP-element group 516: 	 branch_block_stmt_25/bbx_xnph_forx_xbody371_PhiReq/$exit
      -- CP-element group 516: 	 branch_block_stmt_25/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1337/$exit
      -- CP-element group 516: 	 branch_block_stmt_25/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/$exit
      -- CP-element group 516: 	 branch_block_stmt_25/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1341_konst_delay_trans
      -- CP-element group 516: 	 branch_block_stmt_25/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_req
      -- 
    phi_stmt_1337_req_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1337_req_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(516), ack => phi_stmt_1337_req_0); -- 
    -- Element group ct_core_CP_34_elements(516) is a control-delay.
    cp_element_516_delay: control_delay_element  generic map(name => " 516_delay", delay_value => 1)  port map(req => ct_core_CP_34_elements(446), ack => ct_core_CP_34_elements(516), clk => clk, reset =>reset);
    -- CP-element group 517:  transition  input  bypass 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	494 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	519 
    -- CP-element group 517:  members (2) 
      -- CP-element group 517: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/SplitProtocol/Sample/$exit
      -- CP-element group 517: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/SplitProtocol/Sample/ra
      -- 
    ra_3323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1343_inst_ack_0, ack => ct_core_CP_34_elements(517)); -- 
    -- CP-element group 518:  transition  input  bypass 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	494 
    -- CP-element group 518: successors 
    -- CP-element group 518: 	519 
    -- CP-element group 518:  members (2) 
      -- CP-element group 518: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/SplitProtocol/Update/$exit
      -- CP-element group 518: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/SplitProtocol/Update/ca
      -- 
    ca_3328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1343_inst_ack_1, ack => ct_core_CP_34_elements(518)); -- 
    -- CP-element group 519:  join  transition  output  bypass 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	517 
    -- CP-element group 519: 	518 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	520 
    -- CP-element group 519:  members (6) 
      -- CP-element group 519: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/$exit
      -- CP-element group 519: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/$exit
      -- CP-element group 519: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/$exit
      -- CP-element group 519: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/$exit
      -- CP-element group 519: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_sources/type_cast_1343/SplitProtocol/$exit
      -- CP-element group 519: 	 branch_block_stmt_25/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1337/phi_stmt_1337_req
      -- 
    phi_stmt_1337_req_3329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1337_req_3329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(519), ack => phi_stmt_1337_req_1); -- 
    ct_core_cp_element_group_519: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "ct_core_cp_element_group_519"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ct_core_CP_34_elements(517) & ct_core_CP_34_elements(518);
      gj_ct_core_cp_element_group_519 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ct_core_CP_34_elements(519), clk => clk, reset => reset); --
    end block;
    -- CP-element group 520:  merge  transition  place  bypass 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	516 
    -- CP-element group 520: 	519 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	521 
    -- CP-element group 520:  members (2) 
      -- CP-element group 520: 	 branch_block_stmt_25/merge_stmt_1336_PhiReqMerge
      -- CP-element group 520: 	 branch_block_stmt_25/merge_stmt_1336_PhiAck/$entry
      -- 
    ct_core_CP_34_elements(520) <= OrReduce(ct_core_CP_34_elements(516) & ct_core_CP_34_elements(519));
    -- CP-element group 521:  fork  transition  place  input  output  bypass 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	520 
    -- CP-element group 521: successors 
    -- CP-element group 521: 	447 
    -- CP-element group 521: 	448 
    -- CP-element group 521: 	450 
    -- CP-element group 521: 	452 
    -- CP-element group 521: 	454 
    -- CP-element group 521: 	456 
    -- CP-element group 521: 	458 
    -- CP-element group 521: 	460 
    -- CP-element group 521: 	462 
    -- CP-element group 521: 	464 
    -- CP-element group 521: 	466 
    -- CP-element group 521: 	468 
    -- CP-element group 521:  members (53) 
      -- CP-element group 521: 	 branch_block_stmt_25/merge_stmt_1336__exit__
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464__entry__
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_update_start_
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_update_start_
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1418_update_start_
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1378_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1388_update_start_
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1428_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_update_start_
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1368_update_start_
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1408_update_start_
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1398_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_update_start_
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_resized_1
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_scaled_1
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_computed_1
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_resize_1/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_resize_1/$exit
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_resize_1/index_resize_req
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_resize_1/index_resize_ack
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_scale_1/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_scale_1/$exit
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_scale_1/scale_rename_req
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_index_scale_1/scale_rename_ack
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_final_index_sum_regn_update_start
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_final_index_sum_regn_Sample/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_final_index_sum_regn_Sample/req
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_final_index_sum_regn_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/array_obj_ref_1349_final_index_sum_regn_Update/req
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/addr_of_1350_complete/req
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_update_start_
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/word_access_complete/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/word_access_complete/word_0/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/ptr_deref_1354_Update/word_access_complete/word_0/cr
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_update_start_
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_Update/$entry
      -- CP-element group 521: 	 branch_block_stmt_25/assign_stmt_1351_to_assign_stmt_1464/type_cast_1358_Update/cr
      -- CP-element group 521: 	 branch_block_stmt_25/merge_stmt_1336_PhiAck/$exit
      -- CP-element group 521: 	 branch_block_stmt_25/merge_stmt_1336_PhiAck/phi_stmt_1337_ack
      -- 
    phi_stmt_1337_ack_3334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1337_ack_0, ack => ct_core_CP_34_elements(521)); -- 
    cr_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => type_cast_1368_inst_req_1); -- 
    cr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => type_cast_1418_inst_req_1); -- 
    cr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => type_cast_1388_inst_req_1); -- 
    cr_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => type_cast_1378_inst_req_1); -- 
    cr_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => type_cast_1428_inst_req_1); -- 
    cr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => type_cast_1408_inst_req_1); -- 
    cr_2875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => type_cast_1398_inst_req_1); -- 
    req_2735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => array_obj_ref_1349_index_offset_req_0); -- 
    req_2740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => array_obj_ref_1349_index_offset_req_1); -- 
    req_2755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => addr_of_1350_final_reg_req_1); -- 
    cr_2800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => ptr_deref_1354_load_0_req_1); -- 
    cr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ct_core_CP_34_elements(521), ack => type_cast_1358_inst_req_1); -- 
    -- CP-element group 522:  merge  transition  place  bypass 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	444 
    -- CP-element group 522: 	493 
    -- CP-element group 522: successors 
    -- CP-element group 522:  members (16) 
      -- CP-element group 522: 	 $exit
      -- CP-element group 522: 	 branch_block_stmt_25/$exit
      -- CP-element group 522: 	 branch_block_stmt_25/branch_block_stmt_25__exit__
      -- CP-element group 522: 	 branch_block_stmt_25/merge_stmt_1473__exit__
      -- CP-element group 522: 	 branch_block_stmt_25/return__
      -- CP-element group 522: 	 branch_block_stmt_25/merge_stmt_1475__exit__
      -- CP-element group 522: 	 branch_block_stmt_25/merge_stmt_1473_PhiReqMerge
      -- CP-element group 522: 	 branch_block_stmt_25/merge_stmt_1473_PhiAck/$entry
      -- CP-element group 522: 	 branch_block_stmt_25/merge_stmt_1473_PhiAck/$exit
      -- CP-element group 522: 	 branch_block_stmt_25/merge_stmt_1473_PhiAck/dummy
      -- CP-element group 522: 	 branch_block_stmt_25/return___PhiReq/$entry
      -- CP-element group 522: 	 branch_block_stmt_25/return___PhiReq/$exit
      -- CP-element group 522: 	 branch_block_stmt_25/merge_stmt_1475_PhiReqMerge
      -- CP-element group 522: 	 branch_block_stmt_25/merge_stmt_1475_PhiAck/$entry
      -- CP-element group 522: 	 branch_block_stmt_25/merge_stmt_1475_PhiAck/$exit
      -- CP-element group 522: 	 branch_block_stmt_25/merge_stmt_1475_PhiAck/dummy
      -- 
    ct_core_CP_34_elements(522) <= OrReduce(ct_core_CP_34_elements(444) & ct_core_CP_34_elements(493));
    ct_core_do_while_stmt_956_terminator_2396: loop_terminator -- 
      generic map (name => " ct_core_do_while_stmt_956_terminator_2396", max_iterations_in_flight =>15) 
      port map(loop_body_exit => ct_core_CP_34_elements(228),loop_continue => ct_core_CP_34_elements(395),loop_terminate => ct_core_CP_34_elements(394),loop_back => ct_core_CP_34_elements(226),loop_exit => ct_core_CP_34_elements(225),clk => clk, reset => reset); -- 
    phi_stmt_958_phi_seq_1884_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_34_elements(243);
      ct_core_CP_34_elements(246)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_34_elements(246);
      ct_core_CP_34_elements(247)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_34_elements(248);
      ct_core_CP_34_elements(244) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_34_elements(241);
      ct_core_CP_34_elements(250)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_34_elements(252);
      ct_core_CP_34_elements(251)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_34_elements(253);
      ct_core_CP_34_elements(242) <= phi_mux_reqs(1);
      phi_stmt_958_phi_seq_1884 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_958_phi_seq_1884") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_34_elements(233), 
          phi_sample_ack => ct_core_CP_34_elements(239), 
          phi_update_req => ct_core_CP_34_elements(235), 
          phi_update_ack => ct_core_CP_34_elements(240), 
          phi_mux_ack => ct_core_CP_34_elements(245), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_962_phi_seq_1928_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_34_elements(262);
      ct_core_CP_34_elements(265)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_34_elements(265);
      ct_core_CP_34_elements(266)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_34_elements(267);
      ct_core_CP_34_elements(263) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_34_elements(260);
      ct_core_CP_34_elements(269)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_34_elements(271);
      ct_core_CP_34_elements(270)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_34_elements(272);
      ct_core_CP_34_elements(261) <= phi_mux_reqs(1);
      phi_stmt_962_phi_seq_1928 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_962_phi_seq_1928") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_34_elements(256), 
          phi_sample_ack => ct_core_CP_34_elements(257), 
          phi_update_req => ct_core_CP_34_elements(258), 
          phi_update_ack => ct_core_CP_34_elements(259), 
          phi_mux_ack => ct_core_CP_34_elements(264), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_966_phi_seq_1972_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_34_elements(281);
      ct_core_CP_34_elements(284)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_34_elements(284);
      ct_core_CP_34_elements(285)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_34_elements(286);
      ct_core_CP_34_elements(282) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_34_elements(279);
      ct_core_CP_34_elements(288)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_34_elements(290);
      ct_core_CP_34_elements(289)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_34_elements(291);
      ct_core_CP_34_elements(280) <= phi_mux_reqs(1);
      phi_stmt_966_phi_seq_1972 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_966_phi_seq_1972") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_34_elements(275), 
          phi_sample_ack => ct_core_CP_34_elements(276), 
          phi_update_req => ct_core_CP_34_elements(277), 
          phi_update_ack => ct_core_CP_34_elements(278), 
          phi_mux_ack => ct_core_CP_34_elements(283), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_970_phi_seq_2026_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_34_elements(300);
      ct_core_CP_34_elements(303)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_34_elements(305);
      ct_core_CP_34_elements(304)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_34_elements(306);
      ct_core_CP_34_elements(301) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_34_elements(298);
      ct_core_CP_34_elements(307)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_34_elements(309);
      ct_core_CP_34_elements(308)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_34_elements(310);
      ct_core_CP_34_elements(299) <= phi_mux_reqs(1);
      phi_stmt_970_phi_seq_2026 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_970_phi_seq_2026") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_34_elements(294), 
          phi_sample_ack => ct_core_CP_34_elements(295), 
          phi_update_req => ct_core_CP_34_elements(296), 
          phi_update_ack => ct_core_CP_34_elements(297), 
          phi_mux_ack => ct_core_CP_34_elements(302), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_974_phi_seq_2080_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_34_elements(319);
      ct_core_CP_34_elements(322)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_34_elements(324);
      ct_core_CP_34_elements(323)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_34_elements(325);
      ct_core_CP_34_elements(320) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_34_elements(317);
      ct_core_CP_34_elements(326)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_34_elements(328);
      ct_core_CP_34_elements(327)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_34_elements(329);
      ct_core_CP_34_elements(318) <= phi_mux_reqs(1);
      phi_stmt_974_phi_seq_2080 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_974_phi_seq_2080") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_34_elements(313), 
          phi_sample_ack => ct_core_CP_34_elements(314), 
          phi_update_req => ct_core_CP_34_elements(315), 
          phi_update_ack => ct_core_CP_34_elements(316), 
          phi_mux_ack => ct_core_CP_34_elements(321), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_978_phi_seq_2124_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ct_core_CP_34_elements(338);
      ct_core_CP_34_elements(341)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ct_core_CP_34_elements(341);
      ct_core_CP_34_elements(342)<= src_update_reqs(0);
      src_update_acks(0)  <= ct_core_CP_34_elements(343);
      ct_core_CP_34_elements(339) <= phi_mux_reqs(0);
      triggers(1)  <= ct_core_CP_34_elements(336);
      ct_core_CP_34_elements(345)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ct_core_CP_34_elements(347);
      ct_core_CP_34_elements(346)<= src_update_reqs(1);
      src_update_acks(1)  <= ct_core_CP_34_elements(348);
      ct_core_CP_34_elements(337) <= phi_mux_reqs(1);
      phi_stmt_978_phi_seq_2124 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_978_phi_seq_2124") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ct_core_CP_34_elements(332), 
          phi_sample_ack => ct_core_CP_34_elements(333), 
          phi_update_req => ct_core_CP_34_elements(334), 
          phi_update_ack => ct_core_CP_34_elements(335), 
          phi_mux_ack => ct_core_CP_34_elements(340), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1836_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= ct_core_CP_34_elements(229);
        preds(1)  <= ct_core_CP_34_elements(230);
        entry_tmerge_1836 : transition_merge -- 
          generic map(name => " entry_tmerge_1836")
          port map (preds => preds, symbol_out => ct_core_CP_34_elements(231));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal MUX_1118_wire : std_logic_vector(15 downto 0);
    signal MUX_1140_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_1060_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1114_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1136_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1163_wire : std_logic_vector(0 downto 0);
    signal R_indvar469_892_resized : std_logic_vector(13 downto 0);
    signal R_indvar469_892_scaled : std_logic_vector(13 downto 0);
    signal R_indvar476_670_resized : std_logic_vector(9 downto 0);
    signal R_indvar476_670_scaled : std_logic_vector(9 downto 0);
    signal R_indvar489_463_resized : std_logic_vector(13 downto 0);
    signal R_indvar489_463_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1348_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1348_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_1046_1046_delayed_1_0_1052 : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_1142_1142_delayed_1_0_1154 : std_logic_vector(15 downto 0);
    signal add131_491 : std_logic_vector(63 downto 0);
    signal add137_509 : std_logic_vector(63 downto 0);
    signal add143_527 : std_logic_vector(63 downto 0);
    signal add149_545 : std_logic_vector(63 downto 0);
    signal add155_563 : std_logic_vector(63 downto 0);
    signal add161_581 : std_logic_vector(63 downto 0);
    signal add167_599 : std_logic_vector(63 downto 0);
    signal add187_698 : std_logic_vector(63 downto 0);
    signal add193_716 : std_logic_vector(63 downto 0);
    signal add199_734 : std_logic_vector(63 downto 0);
    signal add205_752 : std_logic_vector(63 downto 0);
    signal add211_770 : std_logic_vector(63 downto 0);
    signal add217_788 : std_logic_vector(63 downto 0);
    signal add223_806 : std_logic_vector(63 downto 0);
    signal add_dest_dim0_970 : std_logic_vector(15 downto 0);
    signal add_dest_dim0_init_946 : std_logic_vector(15 downto 0);
    signal add_dest_dim0_init_946_972_buffered : std_logic_vector(15 downto 0);
    signal add_dest_dim1_974 : std_logic_vector(15 downto 0);
    signal add_dest_dim1_init_951 : std_logic_vector(15 downto 0);
    signal add_dest_dim1_init_951_976_buffered : std_logic_vector(15 downto 0);
    signal add_out_1007 : std_logic_vector(15 downto 0);
    signal add_src_978 : std_logic_vector(31 downto 0);
    signal add_src_init_955 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1013_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1013_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1013_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1013_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1013_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1013_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1025_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1349_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1349_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1349_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1349_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1349_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1349_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_464_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_464_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_464_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_464_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_464_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_464_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_671_constant_part_of_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_671_final_offset : std_logic_vector(9 downto 0);
    signal array_obj_ref_671_offset_scale_factor_0 : std_logic_vector(9 downto 0);
    signal array_obj_ref_671_offset_scale_factor_1 : std_logic_vector(9 downto 0);
    signal array_obj_ref_671_resized_base_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_671_root_address : std_logic_vector(9 downto 0);
    signal array_obj_ref_893_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_893_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_893_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_893_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_893_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_893_root_address : std_logic_vector(13 downto 0);
    signal arrayidx227_673 : std_logic_vector(31 downto 0);
    signal arrayidx269_895 : std_logic_vector(31 downto 0);
    signal arrayidx376_1351 : std_logic_vector(31 downto 0);
    signal arrayidx_466 : std_logic_vector(31 downto 0);
    signal call101_229 : std_logic_vector(7 downto 0);
    signal call106_242 : std_logic_vector(7 downto 0);
    signal call10_67 : std_logic_vector(7 downto 0);
    signal call110_254 : std_logic_vector(7 downto 0);
    signal call1124_292 : std_logic_vector(7 downto 0);
    signal call1128_304 : std_logic_vector(7 downto 0);
    signal call115_267 : std_logic_vector(7 downto 0);
    signal call119_279 : std_logic_vector(7 downto 0);
    signal call124_469 : std_logic_vector(7 downto 0);
    signal call128_482 : std_logic_vector(7 downto 0);
    signal call133_317 : std_logic_vector(7 downto 0);
    signal call134_500 : std_logic_vector(7 downto 0);
    signal call140_518 : std_logic_vector(7 downto 0);
    signal call146_536 : std_logic_vector(7 downto 0);
    signal call14_79 : std_logic_vector(7 downto 0);
    signal call152_554 : std_logic_vector(7 downto 0);
    signal call158_572 : std_logic_vector(7 downto 0);
    signal call164_590 : std_logic_vector(7 downto 0);
    signal call180_676 : std_logic_vector(7 downto 0);
    signal call184_689 : std_logic_vector(7 downto 0);
    signal call190_707 : std_logic_vector(7 downto 0);
    signal call196_725 : std_logic_vector(7 downto 0);
    signal call19_92 : std_logic_vector(7 downto 0);
    signal call202_743 : std_logic_vector(7 downto 0);
    signal call208_761 : std_logic_vector(7 downto 0);
    signal call214_779 : std_logic_vector(7 downto 0);
    signal call220_797 : std_logic_vector(7 downto 0);
    signal call233_923 : std_logic_vector(63 downto 0);
    signal call23_104 : std_logic_vector(7 downto 0);
    signal call28_117 : std_logic_vector(7 downto 0);
    signal call297_1170 : std_logic_vector(63 downto 0);
    signal call2_42 : std_logic_vector(7 downto 0);
    signal call32_129 : std_logic_vector(7 downto 0);
    signal call37_142 : std_logic_vector(7 downto 0);
    signal call41_154 : std_logic_vector(7 downto 0);
    signal call46_167 : std_logic_vector(7 downto 0);
    signal call50_179 : std_logic_vector(7 downto 0);
    signal call55_192 : std_logic_vector(7 downto 0);
    signal call5_54 : std_logic_vector(7 downto 0);
    signal call92_204 : std_logic_vector(7 downto 0);
    signal call97_217 : std_logic_vector(7 downto 0);
    signal call_28 : std_logic_vector(7 downto 0);
    signal cmp175463_407 : std_logic_vector(0 downto 0);
    signal cmp264448_836 : std_logic_vector(0 downto 0);
    signal cmp264449_1292 : std_logic_vector(0 downto 0);
    signal cmp467_392 : std_logic_vector(0 downto 0);
    signal cmp_dim0_1063 : std_logic_vector(0 downto 0);
    signal cmp_dim1_1057 : std_logic_vector(0 downto 0);
    signal cmp_dim2_1047 : std_logic_vector(0 downto 0);
    signal continue_flag_1165 : std_logic_vector(0 downto 0);
    signal conv104_233 : std_logic_vector(15 downto 0);
    signal conv107_246 : std_logic_vector(15 downto 0);
    signal conv1125_296 : std_logic_vector(15 downto 0);
    signal conv113_258 : std_logic_vector(15 downto 0);
    signal conv116_271 : std_logic_vector(15 downto 0);
    signal conv11_71 : std_logic_vector(15 downto 0);
    signal conv122_283 : std_logic_vector(15 downto 0);
    signal conv125_473 : std_logic_vector(63 downto 0);
    signal conv130_486 : std_logic_vector(63 downto 0);
    signal conv131_308 : std_logic_vector(15 downto 0);
    signal conv134_321 : std_logic_vector(15 downto 0);
    signal conv136_504 : std_logic_vector(63 downto 0);
    signal conv142_522 : std_logic_vector(63 downto 0);
    signal conv148_540 : std_logic_vector(63 downto 0);
    signal conv154_558 : std_logic_vector(63 downto 0);
    signal conv160_576 : std_logic_vector(63 downto 0);
    signal conv166_594 : std_logic_vector(63 downto 0);
    signal conv17_83 : std_logic_vector(15 downto 0);
    signal conv181_680 : std_logic_vector(63 downto 0);
    signal conv186_693 : std_logic_vector(63 downto 0);
    signal conv192_711 : std_logic_vector(63 downto 0);
    signal conv198_729 : std_logic_vector(63 downto 0);
    signal conv1_33 : std_logic_vector(15 downto 0);
    signal conv204_747 : std_logic_vector(63 downto 0);
    signal conv20_96 : std_logic_vector(15 downto 0);
    signal conv210_765 : std_logic_vector(63 downto 0);
    signal conv216_783 : std_logic_vector(63 downto 0);
    signal conv222_801 : std_logic_vector(63 downto 0);
    signal conv26_108 : std_logic_vector(15 downto 0);
    signal conv276_1176 : std_logic_vector(63 downto 0);
    signal conv298_1181 : std_logic_vector(63 downto 0);
    signal conv29_121 : std_logic_vector(15 downto 0);
    signal conv305_1191 : std_logic_vector(7 downto 0);
    signal conv311_1201 : std_logic_vector(7 downto 0);
    signal conv317_1211 : std_logic_vector(7 downto 0);
    signal conv323_1221 : std_logic_vector(7 downto 0);
    signal conv329_1231 : std_logic_vector(7 downto 0);
    signal conv335_1241 : std_logic_vector(7 downto 0);
    signal conv341_1251 : std_logic_vector(7 downto 0);
    signal conv347_1261 : std_logic_vector(7 downto 0);
    signal conv35_133 : std_logic_vector(15 downto 0);
    signal conv381_1359 : std_logic_vector(7 downto 0);
    signal conv387_1369 : std_logic_vector(7 downto 0);
    signal conv38_146 : std_logic_vector(15 downto 0);
    signal conv393_1379 : std_logic_vector(7 downto 0);
    signal conv399_1389 : std_logic_vector(7 downto 0);
    signal conv3_46 : std_logic_vector(15 downto 0);
    signal conv405_1399 : std_logic_vector(7 downto 0);
    signal conv411_1409 : std_logic_vector(7 downto 0);
    signal conv417_1419 : std_logic_vector(7 downto 0);
    signal conv423_1429 : std_logic_vector(7 downto 0);
    signal conv44_158 : std_logic_vector(15 downto 0);
    signal conv47_171 : std_logic_vector(15 downto 0);
    signal conv53_183 : std_logic_vector(15 downto 0);
    signal conv56_196 : std_logic_vector(15 downto 0);
    signal conv8_58 : std_logic_vector(15 downto 0);
    signal conv95_208 : std_logic_vector(15 downto 0);
    signal conv98_221 : std_logic_vector(15 downto 0);
    signal dim0_end_1159 : std_logic_vector(0 downto 0);
    signal dim2_limit_1039 : std_logic_vector(15 downto 0);
    signal dim2_limit_1039_delayed_1_0_1042 : std_logic_vector(15 downto 0);
    signal exitcond1_1464 : std_logic_vector(0 downto 0);
    signal exitcond22_821 : std_logic_vector(0 downto 0);
    signal exitcond2_614 : std_logic_vector(0 downto 0);
    signal exitcond_911 : std_logic_vector(0 downto 0);
    signal i1_1019 : std_logic_vector(63 downto 0);
    signal iNsTr_111_1321 : std_logic_vector(63 downto 0);
    signal iNsTr_19_436 : std_logic_vector(63 downto 0);
    signal iNsTr_32_643 : std_logic_vector(63 downto 0);
    signal iNsTr_52_865 : std_logic_vector(63 downto 0);
    signal indvar469_881 : std_logic_vector(63 downto 0);
    signal indvar476_659 : std_logic_vector(63 downto 0);
    signal indvar489_452 : std_logic_vector(63 downto 0);
    signal indvar_1337 : std_logic_vector(63 downto 0);
    signal indvarx_xnext470_906 : std_logic_vector(63 downto 0);
    signal indvarx_xnext477_816 : std_logic_vector(63 downto 0);
    signal indvarx_xnext490_609 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1459 : std_logic_vector(63 downto 0);
    signal inp_d0_51 : std_logic_vector(15 downto 0);
    signal inp_d1_76 : std_logic_vector(15 downto 0);
    signal inp_d232_331 : std_logic_vector(31 downto 0);
    signal inp_d2_101 : std_logic_vector(15 downto 0);
    signal input_dim0_958 : std_logic_vector(15 downto 0);
    signal input_dim0_init_928 : std_logic_vector(15 downto 0);
    signal input_dim1_962 : std_logic_vector(15 downto 0);
    signal input_dim1_init_932 : std_logic_vector(15 downto 0);
    signal input_dim2_966 : std_logic_vector(15 downto 0);
    signal input_dim2_init_936 : std_logic_vector(15 downto 0);
    signal input_int1_340 : std_logic_vector(31 downto 0);
    signal input_int_336 : std_logic_vector(15 downto 0);
    signal input_size_345 : std_logic_vector(31 downto 0);
    signal iv1_1015 : std_logic_vector(31 downto 0);
    signal ker_d0_126 : std_logic_vector(15 downto 0);
    signal ker_d1_151 : std_logic_vector(15 downto 0);
    signal ker_d2_176 : std_logic_vector(15 downto 0);
    signal ker_d3_201 : std_logic_vector(15 downto 0);
    signal ker_int1_350 : std_logic_vector(15 downto 0);
    signal ker_int2_355 : std_logic_vector(15 downto 0);
    signal ker_int3_359 : std_logic_vector(31 downto 0);
    signal ker_int4_363 : std_logic_vector(31 downto 0);
    signal kernel_size_368 : std_logic_vector(31 downto 0);
    signal konst_1005_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1037_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1050_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1066_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1071_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1081_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1109_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1131_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1138_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1152_wire_constant : std_logic_vector(15 downto 0);
    signal konst_939_wire_constant : std_logic_vector(15 downto 0);
    signal nao1_992 : std_logic_vector(15 downto 0);
    signal nao2_997 : std_logic_vector(15 downto 0);
    signal nao3_1002 : std_logic_vector(15 downto 0);
    signal nao_987 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim0_1127 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim0_1127_973_buffered : std_logic_vector(15 downto 0);
    signal next_add_dest_dim1_1121 : std_logic_vector(15 downto 0);
    signal next_add_dest_dim1_1121_977_buffered : std_logic_vector(15 downto 0);
    signal next_add_src_1111 : std_logic_vector(31 downto 0);
    signal next_add_src_1111_981_buffered : std_logic_vector(31 downto 0);
    signal next_input_dim0_1149 : std_logic_vector(15 downto 0);
    signal next_input_dim0_1149_961_buffered : std_logic_vector(15 downto 0);
    signal next_input_dim1_1143 : std_logic_vector(15 downto 0);
    signal next_input_dim1_1143_965_buffered : std_logic_vector(15 downto 0);
    signal next_input_dim2_1133 : std_logic_vector(15 downto 0);
    signal next_input_dim2_1133_969_buffered : std_logic_vector(15 downto 0);
    signal nid1_true1_1088 : std_logic_vector(15 downto 0);
    signal nid1_true2_1093 : std_logic_vector(15 downto 0);
    signal nid1_true3_1092_delayed_1_0_1101 : std_logic_vector(15 downto 0);
    signal nid1_true3_1098 : std_logic_vector(15 downto 0);
    signal nid1_true4_1106 : std_logic_vector(15 downto 0);
    signal nid1_true_1083 : std_logic_vector(15 downto 0);
    signal nid2_false1_1078 : std_logic_vector(15 downto 0);
    signal nid2_false_1073 : std_logic_vector(15 downto 0);
    signal nid2_true_1068 : std_logic_vector(15 downto 0);
    signal out_d0_276 : std_logic_vector(15 downto 0);
    signal out_d1_301 : std_logic_vector(15 downto 0);
    signal out_d232_372 : std_logic_vector(31 downto 0);
    signal out_d2_326 : std_logic_vector(15 downto 0);
    signal out_int1_381 : std_logic_vector(31 downto 0);
    signal out_int_377 : std_logic_vector(15 downto 0);
    signal output_size_386 : std_logic_vector(31 downto 0);
    signal ov_1027 : std_logic_vector(31 downto 0);
    signal ov_1028_delayed_6_0_1030 : std_logic_vector(31 downto 0);
    signal pad_941 : std_logic_vector(15 downto 0);
    signal padding_251 : std_logic_vector(15 downto 0);
    signal ptr_deref_1018_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1018_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1018_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1018_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1018_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1032_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1032_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1032_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1032_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1032_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1032_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1354_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1354_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1354_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1354_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1354_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_601_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_601_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_601_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_601_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_601_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_601_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_808_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_808_resized_base_address : std_logic_vector(9 downto 0);
    signal ptr_deref_808_root_address : std_logic_vector(9 downto 0);
    signal ptr_deref_808_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_808_word_address_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_808_word_offset_0 : std_logic_vector(9 downto 0);
    signal ptr_deref_897_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_897_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_897_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_897_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_897_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_897_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_239 : std_logic_vector(15 downto 0);
    signal shl114_264 : std_logic_vector(15 downto 0);
    signal shl123_289 : std_logic_vector(15 downto 0);
    signal shl127_479 : std_logic_vector(63 downto 0);
    signal shl132_314 : std_logic_vector(15 downto 0);
    signal shl133_497 : std_logic_vector(63 downto 0);
    signal shl139_515 : std_logic_vector(63 downto 0);
    signal shl145_533 : std_logic_vector(63 downto 0);
    signal shl151_551 : std_logic_vector(63 downto 0);
    signal shl157_569 : std_logic_vector(63 downto 0);
    signal shl163_587 : std_logic_vector(63 downto 0);
    signal shl183_686 : std_logic_vector(63 downto 0);
    signal shl189_704 : std_logic_vector(63 downto 0);
    signal shl18_89 : std_logic_vector(15 downto 0);
    signal shl195_722 : std_logic_vector(63 downto 0);
    signal shl201_740 : std_logic_vector(63 downto 0);
    signal shl207_758 : std_logic_vector(63 downto 0);
    signal shl213_776 : std_logic_vector(63 downto 0);
    signal shl219_794 : std_logic_vector(63 downto 0);
    signal shl27_114 : std_logic_vector(15 downto 0);
    signal shl36_139 : std_logic_vector(15 downto 0);
    signal shl45_164 : std_logic_vector(15 downto 0);
    signal shl54_189 : std_logic_vector(15 downto 0);
    signal shl96_214 : std_logic_vector(15 downto 0);
    signal shl9_64 : std_logic_vector(15 downto 0);
    signal shl_39 : std_logic_vector(15 downto 0);
    signal shr308_1197 : std_logic_vector(63 downto 0);
    signal shr314_1207 : std_logic_vector(63 downto 0);
    signal shr320_1217 : std_logic_vector(63 downto 0);
    signal shr326_1227 : std_logic_vector(63 downto 0);
    signal shr332_1237 : std_logic_vector(63 downto 0);
    signal shr338_1247 : std_logic_vector(63 downto 0);
    signal shr344_1257 : std_logic_vector(63 downto 0);
    signal shr384_1365 : std_logic_vector(63 downto 0);
    signal shr390_1375 : std_logic_vector(63 downto 0);
    signal shr396_1385 : std_logic_vector(63 downto 0);
    signal shr402_1395 : std_logic_vector(63 downto 0);
    signal shr408_1405 : std_logic_vector(63 downto 0);
    signal shr414_1415 : std_logic_vector(63 downto 0);
    signal shr420_1425 : std_logic_vector(63 downto 0);
    signal stride_226 : std_logic_vector(15 downto 0);
    signal sub_1186 : std_logic_vector(63 downto 0);
    signal tmp377_1355 : std_logic_vector(63 downto 0);
    signal tmp464_1305 : std_logic_vector(31 downto 0);
    signal tmp464x_xop_1317 : std_logic_vector(31 downto 0);
    signal tmp465_1311 : std_logic_vector(0 downto 0);
    signal tmp468_1334 : std_logic_vector(63 downto 0);
    signal tmp476_849 : std_logic_vector(31 downto 0);
    signal tmp476x_xop_861 : std_logic_vector(31 downto 0);
    signal tmp477_855 : std_logic_vector(0 downto 0);
    signal tmp481_878 : std_logic_vector(63 downto 0);
    signal tmp482_627 : std_logic_vector(31 downto 0);
    signal tmp482x_xop_639 : std_logic_vector(31 downto 0);
    signal tmp483_633 : std_logic_vector(0 downto 0);
    signal tmp487_656 : std_logic_vector(63 downto 0);
    signal tmp495_420 : std_logic_vector(31 downto 0);
    signal tmp495x_xop_432 : std_logic_vector(31 downto 0);
    signal tmp496_426 : std_logic_vector(0 downto 0);
    signal tmp500_449 : std_logic_vector(63 downto 0);
    signal type_cast_1012_resized : std_logic_vector(13 downto 0);
    signal type_cast_1012_scaled : std_logic_vector(13 downto 0);
    signal type_cast_1012_wire : std_logic_vector(63 downto 0);
    signal type_cast_1024_resized : std_logic_vector(13 downto 0);
    signal type_cast_1024_scaled : std_logic_vector(13 downto 0);
    signal type_cast_1024_wire : std_logic_vector(63 downto 0);
    signal type_cast_112_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1174_wire : std_logic_vector(63 downto 0);
    signal type_cast_1179_wire : std_logic_vector(63 downto 0);
    signal type_cast_1195_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1205_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1215_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1225_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1235_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1245_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1255_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1290_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1303_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1309_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1315_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1325_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1332_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1341_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1343_wire : std_logic_vector(63 downto 0);
    signal type_cast_1363_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1373_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_137_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1383_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1393_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1403_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1413_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1423_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1457_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_162_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_187_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_212_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_237_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_262_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_287_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_312_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_37_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_390_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_405_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_418_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_424_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_430_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_440_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_447_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_456_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_458_wire : std_logic_vector(63 downto 0);
    signal type_cast_477_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_495_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_531_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_549_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_567_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_585_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_607_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_625_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_62_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_631_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_637_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_647_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_663_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_665_wire : std_logic_vector(63 downto 0);
    signal type_cast_684_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_702_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_720_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_738_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_774_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_792_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_814_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_834_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_847_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_853_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_859_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_869_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_876_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_87_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_885_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_887_wire : std_logic_vector(63 downto 0);
    signal type_cast_899_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_904_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop502_649 : std_logic_vector(63 downto 0);
    signal xx_xop503_442 : std_logic_vector(63 downto 0);
    signal xx_xop513_871 : std_logic_vector(63 downto 0);
    signal xx_xop_1327 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    add_src_init_955 <= "00000000000000000000000000000000";
    array_obj_ref_1013_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1013_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1013_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1013_resized_base_address <= "00000000000000";
    array_obj_ref_1025_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1025_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1025_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1025_resized_base_address <= "00000000000000";
    array_obj_ref_1349_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1349_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1349_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1349_resized_base_address <= "00000000000000";
    array_obj_ref_464_constant_part_of_offset <= "00000000000000";
    array_obj_ref_464_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_464_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_464_resized_base_address <= "00000000000000";
    array_obj_ref_671_constant_part_of_offset <= "0000000000";
    array_obj_ref_671_offset_scale_factor_0 <= "0000000000";
    array_obj_ref_671_offset_scale_factor_1 <= "0000000001";
    array_obj_ref_671_resized_base_address <= "0000000000";
    array_obj_ref_893_constant_part_of_offset <= "00000000000000";
    array_obj_ref_893_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_893_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_893_resized_base_address <= "00000000000000";
    input_dim0_init_928 <= "0000000000000000";
    input_dim1_init_932 <= "0000000000000000";
    input_dim2_init_936 <= "0000000000000000";
    konst_1005_wire_constant <= "0000000000000011";
    konst_1037_wire_constant <= "0000000000001000";
    konst_1050_wire_constant <= "0000000000000001";
    konst_1066_wire_constant <= "0000000000001000";
    konst_1071_wire_constant <= "0000000000000001";
    konst_1081_wire_constant <= "0000000000000001";
    konst_1109_wire_constant <= "00000000000000000000000000000001";
    konst_1131_wire_constant <= "0000000000000000";
    konst_1138_wire_constant <= "0000000000000000";
    konst_1152_wire_constant <= "0000000000000001";
    konst_939_wire_constant <= "0000000000000001";
    ptr_deref_1018_word_offset_0 <= "00000000000000";
    ptr_deref_1032_word_offset_0 <= "00000000000000";
    ptr_deref_1354_word_offset_0 <= "00000000000000";
    ptr_deref_601_word_offset_0 <= "00000000000000";
    ptr_deref_808_word_offset_0 <= "0000000000";
    ptr_deref_897_word_offset_0 <= "00000000000000";
    type_cast_112_wire_constant <= "0000000000001000";
    type_cast_1195_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1205_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1215_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1225_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1235_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1245_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1255_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1290_wire_constant <= "00000000000000000000000000000111";
    type_cast_1303_wire_constant <= "00000000000000000000000000000011";
    type_cast_1309_wire_constant <= "00000000000000000000000000000001";
    type_cast_1315_wire_constant <= "11111111111111111111111111111111";
    type_cast_1325_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1332_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1341_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1363_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1373_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_137_wire_constant <= "0000000000001000";
    type_cast_1383_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1393_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1403_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1413_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1423_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1457_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_162_wire_constant <= "0000000000001000";
    type_cast_187_wire_constant <= "0000000000001000";
    type_cast_212_wire_constant <= "0000000000001000";
    type_cast_237_wire_constant <= "0000000000001000";
    type_cast_262_wire_constant <= "0000000000001000";
    type_cast_287_wire_constant <= "0000000000001000";
    type_cast_312_wire_constant <= "0000000000001000";
    type_cast_37_wire_constant <= "0000000000001000";
    type_cast_390_wire_constant <= "00000000000000000000000000000111";
    type_cast_405_wire_constant <= "00000000000000000000000000000111";
    type_cast_418_wire_constant <= "00000000000000000000000000000011";
    type_cast_424_wire_constant <= "00000000000000000000000000000001";
    type_cast_430_wire_constant <= "11111111111111111111111111111111";
    type_cast_440_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_447_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_456_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_477_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_495_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_513_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_531_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_549_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_567_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_585_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_607_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_625_wire_constant <= "00000000000000000000000000000011";
    type_cast_62_wire_constant <= "0000000000001000";
    type_cast_631_wire_constant <= "00000000000000000000000000000001";
    type_cast_637_wire_constant <= "11111111111111111111111111111111";
    type_cast_647_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_654_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_663_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_684_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_702_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_720_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_738_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_756_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_774_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_792_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_814_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_834_wire_constant <= "00000000000000000000000000000011";
    type_cast_847_wire_constant <= "00000000000000000000000000000011";
    type_cast_853_wire_constant <= "00000000000000000000000000000001";
    type_cast_859_wire_constant <= "11111111111111111111111111111111";
    type_cast_869_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_876_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_87_wire_constant <= "0000000000001000";
    type_cast_885_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_899_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_904_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1337: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1341_wire_constant & type_cast_1343_wire;
      req <= phi_stmt_1337_req_0 & phi_stmt_1337_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1337",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1337_ack_0,
          idata => idata,
          odata => indvar_1337,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1337
    phi_stmt_452: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_456_wire_constant & type_cast_458_wire;
      req <= phi_stmt_452_req_0 & phi_stmt_452_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_452",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_452_ack_0,
          idata => idata,
          odata => indvar489_452,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_452
    phi_stmt_659: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_663_wire_constant & type_cast_665_wire;
      req <= phi_stmt_659_req_0 & phi_stmt_659_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_659",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_659_ack_0,
          idata => idata,
          odata => indvar476_659,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_659
    phi_stmt_881: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_885_wire_constant & type_cast_887_wire;
      req <= phi_stmt_881_req_0 & phi_stmt_881_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_881",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_881_ack_0,
          idata => idata,
          odata => indvar469_881,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_881
    phi_stmt_958: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim0_init_928 & next_input_dim0_1149_961_buffered;
      req <= phi_stmt_958_req_0 & phi_stmt_958_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_958",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_958_ack_0,
          idata => idata,
          odata => input_dim0_958,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_958
    phi_stmt_962: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim1_init_932 & next_input_dim1_1143_965_buffered;
      req <= phi_stmt_962_req_0 & phi_stmt_962_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_962",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_962_ack_0,
          idata => idata,
          odata => input_dim1_962,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_962
    phi_stmt_966: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= input_dim2_init_936 & next_input_dim2_1133_969_buffered;
      req <= phi_stmt_966_req_0 & phi_stmt_966_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_966",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_966_ack_0,
          idata => idata,
          odata => input_dim2_966,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_966
    phi_stmt_970: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_dest_dim0_init_946_972_buffered & next_add_dest_dim0_1127_973_buffered;
      req <= phi_stmt_970_req_0 & phi_stmt_970_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_970",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_970_ack_0,
          idata => idata,
          odata => add_dest_dim0_970,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_970
    phi_stmt_974: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_dest_dim1_init_951_976_buffered & next_add_dest_dim1_1121_977_buffered;
      req <= phi_stmt_974_req_0 & phi_stmt_974_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_974",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_974_ack_0,
          idata => idata,
          odata => add_dest_dim1_974,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_974
    phi_stmt_978: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_src_init_955 & next_add_src_1111_981_buffered;
      req <= phi_stmt_978_req_0 & phi_stmt_978_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_978",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_978_ack_0,
          idata => idata,
          odata => add_src_978,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_978
    -- flow-through select operator MUX_1118_inst
    MUX_1118_wire <= nid1_true4_1106 when (cmp_dim1_1057(0) /=  '0') else nid2_false1_1078;
    -- flow-through select operator MUX_1120_inst
    next_add_dest_dim1_1121 <= MUX_1118_wire when (NOT_u1_u1_1114_wire(0) /=  '0') else add_dest_dim1_974;
    -- flow-through select operator MUX_1126_inst
    next_add_dest_dim0_1127 <= nid1_true1_1088 when (cmp_dim0_1063(0) /=  '0') else add_dest_dim0_970;
    -- flow-through select operator MUX_1132_inst
    next_input_dim2_1133 <= nid2_true_1068 when (cmp_dim2_1047(0) /=  '0') else konst_1131_wire_constant;
    -- flow-through select operator MUX_1140_inst
    MUX_1140_wire <= konst_1138_wire_constant when (cmp_dim1_1057(0) /=  '0') else nid2_false_1073;
    -- flow-through select operator MUX_1142_inst
    next_input_dim1_1143 <= MUX_1140_wire when (NOT_u1_u1_1136_wire(0) /=  '0') else input_dim1_962;
    -- flow-through select operator MUX_1148_inst
    next_input_dim0_1149 <= nid1_true_1083 when (cmp_dim0_1063(0) /=  '0') else input_dim0_958;
    -- flow-through select operator MUX_1333_inst
    tmp468_1334 <= xx_xop_1327 when (tmp465_1311(0) /=  '0') else type_cast_1332_wire_constant;
    -- flow-through select operator MUX_448_inst
    tmp500_449 <= xx_xop503_442 when (tmp496_426(0) /=  '0') else type_cast_447_wire_constant;
    -- flow-through select operator MUX_655_inst
    tmp487_656 <= xx_xop502_649 when (tmp483_633(0) /=  '0') else type_cast_654_wire_constant;
    -- flow-through select operator MUX_877_inst
    tmp481_878 <= xx_xop513_871 when (tmp477_855(0) /=  '0') else type_cast_876_wire_constant;
    W_dim2_limit_1039_delayed_1_0_1040_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_dim2_limit_1039_delayed_1_0_1040_inst_req_0;
      W_dim2_limit_1039_delayed_1_0_1040_inst_ack_0<= wack(0);
      rreq(0) <= W_dim2_limit_1039_delayed_1_0_1040_inst_req_1;
      W_dim2_limit_1039_delayed_1_0_1040_inst_ack_1<= rack(0);
      W_dim2_limit_1039_delayed_1_0_1040_inst : InterlockBuffer generic map ( -- 
        name => "W_dim2_limit_1039_delayed_1_0_1040_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => dim2_limit_1039,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => dim2_limit_1039_delayed_1_0_1042,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_nid1_true3_1092_delayed_1_0_1099_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_nid1_true3_1092_delayed_1_0_1099_inst_req_0;
      W_nid1_true3_1092_delayed_1_0_1099_inst_ack_0<= wack(0);
      rreq(0) <= W_nid1_true3_1092_delayed_1_0_1099_inst_req_1;
      W_nid1_true3_1092_delayed_1_0_1099_inst_ack_1<= rack(0);
      W_nid1_true3_1092_delayed_1_0_1099_inst : InterlockBuffer generic map ( -- 
        name => "W_nid1_true3_1092_delayed_1_0_1099_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nid1_true3_1098,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nid1_true3_1092_delayed_1_0_1101,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ov_1028_delayed_6_0_1028_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ov_1028_delayed_6_0_1028_inst_req_0;
      W_ov_1028_delayed_6_0_1028_inst_ack_0<= wack(0);
      rreq(0) <= W_ov_1028_delayed_6_0_1028_inst_req_1;
      W_ov_1028_delayed_6_0_1028_inst_ack_1<= rack(0);
      W_ov_1028_delayed_6_0_1028_inst : InterlockBuffer generic map ( -- 
        name => "W_ov_1028_delayed_6_0_1028_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ov_1027,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ov_1028_delayed_6_0_1030,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    add_dest_dim0_init_946_972_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= add_dest_dim0_init_946_972_buf_req_0;
      add_dest_dim0_init_946_972_buf_ack_0<= wack(0);
      rreq(0) <= add_dest_dim0_init_946_972_buf_req_1;
      add_dest_dim0_init_946_972_buf_ack_1<= rack(0);
      add_dest_dim0_init_946_972_buf : InterlockBuffer generic map ( -- 
        name => "add_dest_dim0_init_946_972_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim0_init_946,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim0_init_946_972_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    add_dest_dim1_init_951_976_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= add_dest_dim1_init_951_976_buf_req_0;
      add_dest_dim1_init_951_976_buf_ack_0<= wack(0);
      rreq(0) <= add_dest_dim1_init_951_976_buf_req_1;
      add_dest_dim1_init_951_976_buf_ack_1<= rack(0);
      add_dest_dim1_init_951_976_buf : InterlockBuffer generic map ( -- 
        name => "add_dest_dim1_init_951_976_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_dest_dim1_init_951,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_dest_dim1_init_951_976_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1014_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1014_final_reg_req_0;
      addr_of_1014_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1014_final_reg_req_1;
      addr_of_1014_final_reg_ack_1<= rack(0);
      addr_of_1014_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1014_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1013_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iv1_1015,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1026_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1026_final_reg_req_0;
      addr_of_1026_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1026_final_reg_req_1;
      addr_of_1026_final_reg_ack_1<= rack(0);
      addr_of_1026_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1026_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1025_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ov_1027,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1350_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1350_final_reg_req_0;
      addr_of_1350_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1350_final_reg_req_1;
      addr_of_1350_final_reg_ack_1<= rack(0);
      addr_of_1350_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1350_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1349_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx376_1351,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_465_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_465_final_reg_req_0;
      addr_of_465_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_465_final_reg_req_1;
      addr_of_465_final_reg_ack_1<= rack(0);
      addr_of_465_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_465_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_464_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_466,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_672_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_672_final_reg_req_0;
      addr_of_672_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_672_final_reg_req_1;
      addr_of_672_final_reg_ack_1<= rack(0);
      addr_of_672_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_672_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 10,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_671_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx227_673,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_894_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_894_final_reg_req_0;
      addr_of_894_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_894_final_reg_req_1;
      addr_of_894_final_reg_ack_1<= rack(0);
      addr_of_894_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_894_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_893_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_895,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_dest_dim0_1127_973_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_dest_dim0_1127_973_buf_req_0;
      next_add_dest_dim0_1127_973_buf_ack_0<= wack(0);
      rreq(0) <= next_add_dest_dim0_1127_973_buf_req_1;
      next_add_dest_dim0_1127_973_buf_ack_1<= rack(0);
      next_add_dest_dim0_1127_973_buf : InterlockBuffer generic map ( -- 
        name => "next_add_dest_dim0_1127_973_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_dest_dim0_1127,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_dest_dim0_1127_973_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_dest_dim1_1121_977_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_dest_dim1_1121_977_buf_req_0;
      next_add_dest_dim1_1121_977_buf_ack_0<= wack(0);
      rreq(0) <= next_add_dest_dim1_1121_977_buf_req_1;
      next_add_dest_dim1_1121_977_buf_ack_1<= rack(0);
      next_add_dest_dim1_1121_977_buf : InterlockBuffer generic map ( -- 
        name => "next_add_dest_dim1_1121_977_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_dest_dim1_1121,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_dest_dim1_1121_977_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_src_1111_981_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_src_1111_981_buf_req_0;
      next_add_src_1111_981_buf_ack_0<= wack(0);
      rreq(0) <= next_add_src_1111_981_buf_req_1;
      next_add_src_1111_981_buf_ack_1<= rack(0);
      next_add_src_1111_981_buf : InterlockBuffer generic map ( -- 
        name => "next_add_src_1111_981_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_src_1111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_src_1111_981_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim0_1149_961_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim0_1149_961_buf_req_0;
      next_input_dim0_1149_961_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim0_1149_961_buf_req_1;
      next_input_dim0_1149_961_buf_ack_1<= rack(0);
      next_input_dim0_1149_961_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim0_1149_961_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim0_1149,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim0_1149_961_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim1_1143_965_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim1_1143_965_buf_req_0;
      next_input_dim1_1143_965_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim1_1143_965_buf_req_1;
      next_input_dim1_1143_965_buf_ack_1<= rack(0);
      next_input_dim1_1143_965_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim1_1143_965_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim1_1143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim1_1143_965_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_input_dim2_1133_969_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_input_dim2_1133_969_buf_req_0;
      next_input_dim2_1133_969_buf_ack_0<= wack(0);
      rreq(0) <= next_input_dim2_1133_969_buf_req_1;
      next_input_dim2_1133_969_buf_ack_1<= rack(0);
      next_input_dim2_1133_969_buf : InterlockBuffer generic map ( -- 
        name => "next_input_dim2_1133_969_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_input_dim2_1133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_input_dim2_1133_969_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1012_inst
    process(add_src_978) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_src_978(31 downto 0);
      type_cast_1012_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1024_inst
    process(add_out_1007) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := add_out_1007(15 downto 0);
      type_cast_1024_wire <= tmp_var; -- 
    end process;
    type_cast_107_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_107_inst_req_0;
      type_cast_107_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_107_inst_req_1;
      type_cast_107_inst_ack_1<= rack(0);
      type_cast_107_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_107_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_104,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_108,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1175_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1175_inst_req_0;
      type_cast_1175_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1175_inst_req_1;
      type_cast_1175_inst_ack_1<= rack(0);
      type_cast_1175_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1175_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1174_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_1176,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1180_inst_req_0;
      type_cast_1180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1180_inst_req_1;
      type_cast_1180_inst_ack_1<= rack(0);
      type_cast_1180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1179_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv298_1181,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1190_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1190_inst_req_0;
      type_cast_1190_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1190_inst_req_1;
      type_cast_1190_inst_ack_1<= rack(0);
      type_cast_1190_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1190_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1191,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1200_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1200_inst_req_0;
      type_cast_1200_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1200_inst_req_1;
      type_cast_1200_inst_ack_1<= rack(0);
      type_cast_1200_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1200_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr308_1197,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv311_1201,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_120_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_120_inst_req_0;
      type_cast_120_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_120_inst_req_1;
      type_cast_120_inst_ack_1<= rack(0);
      type_cast_120_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_120_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1210_inst_req_0;
      type_cast_1210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1210_inst_req_1;
      type_cast_1210_inst_ack_1<= rack(0);
      type_cast_1210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr314_1207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv317_1211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1220_inst_req_0;
      type_cast_1220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1220_inst_req_1;
      type_cast_1220_inst_ack_1<= rack(0);
      type_cast_1220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr320_1217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv323_1221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1230_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1230_inst_req_0;
      type_cast_1230_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1230_inst_req_1;
      type_cast_1230_inst_ack_1<= rack(0);
      type_cast_1230_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1230_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr326_1227,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv329_1231,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1240_inst_req_0;
      type_cast_1240_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1240_inst_req_1;
      type_cast_1240_inst_ack_1<= rack(0);
      type_cast_1240_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1240_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr332_1237,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv335_1241,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1250_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1250_inst_req_0;
      type_cast_1250_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1250_inst_req_1;
      type_cast_1250_inst_ack_1<= rack(0);
      type_cast_1250_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1250_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1251,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1260_inst_req_0;
      type_cast_1260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1260_inst_req_1;
      type_cast_1260_inst_ack_1<= rack(0);
      type_cast_1260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr344_1257,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv347_1261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1320_inst_req_0;
      type_cast_1320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1320_inst_req_1;
      type_cast_1320_inst_ack_1<= rack(0);
      type_cast_1320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp464x_xop_1317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_111_1321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_132_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_132_inst_req_0;
      type_cast_132_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_132_inst_req_1;
      type_cast_132_inst_ack_1<= rack(0);
      type_cast_132_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_132_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_133,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1343_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1343_inst_req_0;
      type_cast_1343_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1343_inst_req_1;
      type_cast_1343_inst_ack_1<= rack(0);
      type_cast_1343_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1343_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1459,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1343_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1358_inst_req_0;
      type_cast_1358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1358_inst_req_1;
      type_cast_1358_inst_ack_1<= rack(0);
      type_cast_1358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp377_1355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv381_1359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1368_inst_req_0;
      type_cast_1368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1368_inst_req_1;
      type_cast_1368_inst_ack_1<= rack(0);
      type_cast_1368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr384_1365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv387_1369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1378_inst_req_0;
      type_cast_1378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1378_inst_req_1;
      type_cast_1378_inst_ack_1<= rack(0);
      type_cast_1378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr390_1375,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv393_1379,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1388_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1388_inst_req_0;
      type_cast_1388_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1388_inst_req_1;
      type_cast_1388_inst_ack_1<= rack(0);
      type_cast_1388_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1388_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr396_1385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv399_1389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1398_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1398_inst_req_0;
      type_cast_1398_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1398_inst_req_1;
      type_cast_1398_inst_ack_1<= rack(0);
      type_cast_1398_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1398_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr402_1395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv405_1399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1408_inst_req_0;
      type_cast_1408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1408_inst_req_1;
      type_cast_1408_inst_ack_1<= rack(0);
      type_cast_1408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1408_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr408_1405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv411_1409,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1418_inst_req_0;
      type_cast_1418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1418_inst_req_1;
      type_cast_1418_inst_ack_1<= rack(0);
      type_cast_1418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr414_1415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv417_1419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1428_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1428_inst_req_0;
      type_cast_1428_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1428_inst_req_1;
      type_cast_1428_inst_ack_1<= rack(0);
      type_cast_1428_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1428_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr420_1425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv423_1429,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_145_inst_req_0;
      type_cast_145_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_145_inst_req_1;
      type_cast_145_inst_ack_1<= rack(0);
      type_cast_145_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_145_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_146,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_157_inst_req_0;
      type_cast_157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_157_inst_req_1;
      type_cast_157_inst_ack_1<= rack(0);
      type_cast_157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_170_inst_req_0;
      type_cast_170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_170_inst_req_1;
      type_cast_170_inst_ack_1<= rack(0);
      type_cast_170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_182_inst_req_0;
      type_cast_182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_182_inst_req_1;
      type_cast_182_inst_ack_1<= rack(0);
      type_cast_182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_195_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_195_inst_req_0;
      type_cast_195_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_195_inst_req_1;
      type_cast_195_inst_ack_1<= rack(0);
      type_cast_195_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_195_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_196,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_207_inst_req_0;
      type_cast_207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_207_inst_req_1;
      type_cast_207_inst_ack_1<= rack(0);
      type_cast_207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_220_inst_req_0;
      type_cast_220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_220_inst_req_1;
      type_cast_220_inst_ack_1<= rack(0);
      type_cast_220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_232_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_232_inst_req_0;
      type_cast_232_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_232_inst_req_1;
      type_cast_232_inst_ack_1<= rack(0);
      type_cast_232_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_232_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_229,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_233,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_245_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_245_inst_req_0;
      type_cast_245_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_245_inst_req_1;
      type_cast_245_inst_ack_1<= rack(0);
      type_cast_245_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_245_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_242,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_246,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_257_inst_req_0;
      type_cast_257_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_257_inst_req_1;
      type_cast_257_inst_ack_1<= rack(0);
      type_cast_257_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_257_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_258,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_270_inst_req_0;
      type_cast_270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_270_inst_req_1;
      type_cast_270_inst_ack_1<= rack(0);
      type_cast_270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_270_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_267,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_282_inst_req_0;
      type_cast_282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_282_inst_req_1;
      type_cast_282_inst_ack_1<= rack(0);
      type_cast_282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_279,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_283,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_295_inst_req_0;
      type_cast_295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_295_inst_req_1;
      type_cast_295_inst_ack_1<= rack(0);
      type_cast_295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1124_292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1125_296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_307_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_307_inst_req_0;
      type_cast_307_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_307_inst_req_1;
      type_cast_307_inst_ack_1<= rack(0);
      type_cast_307_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_307_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1128_304,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_308,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_320_inst_req_0;
      type_cast_320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_320_inst_req_1;
      type_cast_320_inst_ack_1<= rack(0);
      type_cast_320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_32_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_32_inst_req_0;
      type_cast_32_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_32_inst_req_1;
      type_cast_32_inst_ack_1<= rack(0);
      type_cast_32_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_32_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_28,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_33,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_330_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_330_inst_req_0;
      type_cast_330_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_330_inst_req_1;
      type_cast_330_inst_ack_1<= rack(0);
      type_cast_330_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_330_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inp_d2_101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inp_d232_331,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_339_inst_req_0;
      type_cast_339_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_339_inst_req_1;
      type_cast_339_inst_ack_1<= rack(0);
      type_cast_339_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_int_336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_int1_340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_358_inst_req_0;
      type_cast_358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_358_inst_req_1;
      type_cast_358_inst_ack_1<= rack(0);
      type_cast_358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ker_int1_350,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ker_int3_359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_362_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_362_inst_req_0;
      type_cast_362_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_362_inst_req_1;
      type_cast_362_inst_ack_1<= rack(0);
      type_cast_362_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_362_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ker_int2_355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ker_int4_363,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_371_inst_req_0;
      type_cast_371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_371_inst_req_1;
      type_cast_371_inst_ack_1<= rack(0);
      type_cast_371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inp_d2_101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => out_d232_372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_380_inst_req_0;
      type_cast_380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_380_inst_req_1;
      type_cast_380_inst_ack_1<= rack(0);
      type_cast_380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => out_int_377,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => out_int1_381,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_435_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_435_inst_req_0;
      type_cast_435_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_435_inst_req_1;
      type_cast_435_inst_ack_1<= rack(0);
      type_cast_435_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_435_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp495x_xop_432,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_19_436,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_458_inst_req_0;
      type_cast_458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_458_inst_req_1;
      type_cast_458_inst_ack_1<= rack(0);
      type_cast_458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_458_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext490_609,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_458_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_45_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_45_inst_req_0;
      type_cast_45_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_45_inst_req_1;
      type_cast_45_inst_ack_1<= rack(0);
      type_cast_45_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_45_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_42,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_46,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_472_inst_req_0;
      type_cast_472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_472_inst_req_1;
      type_cast_472_inst_ack_1<= rack(0);
      type_cast_472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_469,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_485_inst_req_0;
      type_cast_485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_485_inst_req_1;
      type_cast_485_inst_ack_1<= rack(0);
      type_cast_485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_503_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_503_inst_req_0;
      type_cast_503_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_503_inst_req_1;
      type_cast_503_inst_ack_1<= rack(0);
      type_cast_503_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_503_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call134_500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv136_504,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_521_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_521_inst_req_0;
      type_cast_521_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_521_inst_req_1;
      type_cast_521_inst_ack_1<= rack(0);
      type_cast_521_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_521_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call140_518,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv142_522,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_539_inst_req_0;
      type_cast_539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_539_inst_req_1;
      type_cast_539_inst_ack_1<= rack(0);
      type_cast_539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call146_536,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv148_540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_557_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_557_inst_req_0;
      type_cast_557_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_557_inst_req_1;
      type_cast_557_inst_ack_1<= rack(0);
      type_cast_557_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_557_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call152_554,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_558,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_575_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_575_inst_req_0;
      type_cast_575_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_575_inst_req_1;
      type_cast_575_inst_ack_1<= rack(0);
      type_cast_575_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_575_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call158_572,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv160_576,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_57_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_57_inst_req_0;
      type_cast_57_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_57_inst_req_1;
      type_cast_57_inst_ack_1<= rack(0);
      type_cast_57_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_57_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_54,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_58,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_593_inst_req_0;
      type_cast_593_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_593_inst_req_1;
      type_cast_593_inst_ack_1<= rack(0);
      type_cast_593_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_593_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_590,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv166_594,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_642_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_642_inst_req_0;
      type_cast_642_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_642_inst_req_1;
      type_cast_642_inst_ack_1<= rack(0);
      type_cast_642_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_642_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp482x_xop_639,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_32_643,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_665_inst_req_0;
      type_cast_665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_665_inst_req_1;
      type_cast_665_inst_ack_1<= rack(0);
      type_cast_665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_665_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext477_816,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_665_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_679_inst_req_0;
      type_cast_679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_679_inst_req_1;
      type_cast_679_inst_ack_1<= rack(0);
      type_cast_679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_679_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_676,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv181_680,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_692_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_692_inst_req_0;
      type_cast_692_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_692_inst_req_1;
      type_cast_692_inst_ack_1<= rack(0);
      type_cast_692_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_692_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call184_689,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv186_693,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_70_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_70_inst_req_0;
      type_cast_70_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_70_inst_req_1;
      type_cast_70_inst_ack_1<= rack(0);
      type_cast_70_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_70_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_67,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_71,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_710_inst_req_0;
      type_cast_710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_710_inst_req_1;
      type_cast_710_inst_ack_1<= rack(0);
      type_cast_710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call190_707,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv192_711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_728_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_728_inst_req_0;
      type_cast_728_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_728_inst_req_1;
      type_cast_728_inst_ack_1<= rack(0);
      type_cast_728_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_728_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call196_725,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv198_729,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_746_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_746_inst_req_0;
      type_cast_746_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_746_inst_req_1;
      type_cast_746_inst_ack_1<= rack(0);
      type_cast_746_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_746_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call202_743,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv204_747,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_764_inst_req_0;
      type_cast_764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_764_inst_req_1;
      type_cast_764_inst_ack_1<= rack(0);
      type_cast_764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call208_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv210_765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_782_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_782_inst_req_0;
      type_cast_782_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_782_inst_req_1;
      type_cast_782_inst_ack_1<= rack(0);
      type_cast_782_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_782_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call214_779,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv216_783,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_800_inst_req_0;
      type_cast_800_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_800_inst_req_1;
      type_cast_800_inst_ack_1<= rack(0);
      type_cast_800_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_800_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call220_797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv222_801,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_82_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_82_inst_req_0;
      type_cast_82_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_82_inst_req_1;
      type_cast_82_inst_ack_1<= rack(0);
      type_cast_82_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_82_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_79,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_83,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_864_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_864_inst_req_0;
      type_cast_864_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_864_inst_req_1;
      type_cast_864_inst_ack_1<= rack(0);
      type_cast_864_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_864_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp476x_xop_861,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_52_865,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_887_inst_req_0;
      type_cast_887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_887_inst_req_1;
      type_cast_887_inst_ack_1<= rack(0);
      type_cast_887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext470_906,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_887_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_95_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_95_inst_req_0;
      type_cast_95_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_95_inst_req_1;
      type_cast_95_inst_ack_1<= rack(0);
      type_cast_95_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_95_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_92,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_96,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1013_index_1_rename
    process(type_cast_1012_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1012_resized;
      ov(13 downto 0) := iv;
      type_cast_1012_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1013_index_1_resize
    process(type_cast_1012_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1012_wire;
      ov := iv(13 downto 0);
      type_cast_1012_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1013_root_address_inst
    process(array_obj_ref_1013_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1013_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1013_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1025_index_1_rename
    process(type_cast_1024_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1024_resized;
      ov(13 downto 0) := iv;
      type_cast_1024_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1025_index_1_resize
    process(type_cast_1024_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1024_wire;
      ov := iv(13 downto 0);
      type_cast_1024_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1025_root_address_inst
    process(array_obj_ref_1025_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1025_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1025_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1349_index_1_rename
    process(R_indvar_1348_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1348_resized;
      ov(13 downto 0) := iv;
      R_indvar_1348_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1349_index_1_resize
    process(indvar_1337) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1337;
      ov := iv(13 downto 0);
      R_indvar_1348_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1349_root_address_inst
    process(array_obj_ref_1349_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1349_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1349_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_464_index_1_rename
    process(R_indvar489_463_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar489_463_resized;
      ov(13 downto 0) := iv;
      R_indvar489_463_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_464_index_1_resize
    process(indvar489_452) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar489_452;
      ov := iv(13 downto 0);
      R_indvar489_463_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_464_root_address_inst
    process(array_obj_ref_464_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_464_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_464_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_671_index_1_rename
    process(R_indvar476_670_resized) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar476_670_resized;
      ov(9 downto 0) := iv;
      R_indvar476_670_scaled <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_671_index_1_resize
    process(indvar476_659) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar476_659;
      ov := iv(9 downto 0);
      R_indvar476_670_resized <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_671_root_address_inst
    process(array_obj_ref_671_final_offset) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_671_final_offset;
      ov(9 downto 0) := iv;
      array_obj_ref_671_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_893_index_1_rename
    process(R_indvar469_892_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar469_892_resized;
      ov(13 downto 0) := iv;
      R_indvar469_892_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_893_index_1_resize
    process(indvar469_881) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar469_881;
      ov := iv(13 downto 0);
      R_indvar469_892_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_893_root_address_inst
    process(array_obj_ref_893_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_893_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_893_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1018_addr_0
    process(ptr_deref_1018_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1018_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1018_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1018_base_resize
    process(iv1_1015) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iv1_1015;
      ov := iv(13 downto 0);
      ptr_deref_1018_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1018_gather_scatter
    process(ptr_deref_1018_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1018_data_0;
      ov(63 downto 0) := iv;
      i1_1019 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1018_root_address_inst
    process(ptr_deref_1018_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1018_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1018_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1032_addr_0
    process(ptr_deref_1032_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1032_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1032_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1032_base_resize
    process(ov_1028_delayed_6_0_1030) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ov_1028_delayed_6_0_1030;
      ov := iv(13 downto 0);
      ptr_deref_1032_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1032_gather_scatter
    process(i1_1019) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := i1_1019;
      ov(63 downto 0) := iv;
      ptr_deref_1032_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1032_root_address_inst
    process(ptr_deref_1032_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1032_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1032_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1354_addr_0
    process(ptr_deref_1354_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1354_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1354_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1354_base_resize
    process(arrayidx376_1351) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx376_1351;
      ov := iv(13 downto 0);
      ptr_deref_1354_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1354_gather_scatter
    process(ptr_deref_1354_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1354_data_0;
      ov(63 downto 0) := iv;
      tmp377_1355 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1354_root_address_inst
    process(ptr_deref_1354_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1354_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1354_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_601_addr_0
    process(ptr_deref_601_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_601_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_601_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_601_base_resize
    process(arrayidx_466) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_466;
      ov := iv(13 downto 0);
      ptr_deref_601_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_601_gather_scatter
    process(add167_599) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add167_599;
      ov(63 downto 0) := iv;
      ptr_deref_601_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_601_root_address_inst
    process(ptr_deref_601_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_601_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_601_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_808_addr_0
    process(ptr_deref_808_root_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_808_root_address;
      ov(9 downto 0) := iv;
      ptr_deref_808_word_address_0 <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_808_base_resize
    process(arrayidx227_673) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx227_673;
      ov := iv(9 downto 0);
      ptr_deref_808_resized_base_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_808_gather_scatter
    process(add223_806) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add223_806;
      ov(63 downto 0) := iv;
      ptr_deref_808_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_808_root_address_inst
    process(ptr_deref_808_resized_base_address) --
      variable iv : std_logic_vector(9 downto 0);
      variable ov : std_logic_vector(9 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_808_resized_base_address;
      ov(9 downto 0) := iv;
      ptr_deref_808_root_address <= ov(9 downto 0);
      --
    end process;
    -- equivalence ptr_deref_897_addr_0
    process(ptr_deref_897_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_897_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_897_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_897_base_resize
    process(arrayidx269_895) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_895;
      ov := iv(13 downto 0);
      ptr_deref_897_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_897_gather_scatter
    process(type_cast_899_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_899_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_897_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_897_root_address_inst
    process(ptr_deref_897_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_897_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_897_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_956_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_1165;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_956_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_956_branch_req_0,
          ack0 => do_while_stmt_956_branch_ack_0,
          ack1 => do_while_stmt_956_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1293_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264449_1292;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1293_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1293_branch_req_0,
          ack0 => if_stmt_1293_branch_ack_0,
          ack1 => if_stmt_1293_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1465_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1464;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1465_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1465_branch_req_0,
          ack0 => if_stmt_1465_branch_ack_0,
          ack1 => if_stmt_1465_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_393_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp467_392;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_393_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_393_branch_req_0,
          ack0 => if_stmt_393_branch_ack_0,
          ack1 => if_stmt_393_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_408_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp175463_407;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_408_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_408_branch_req_0,
          ack0 => if_stmt_408_branch_ack_0,
          ack1 => if_stmt_408_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_615_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_614;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_615_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_615_branch_req_0,
          ack0 => if_stmt_615_branch_ack_0,
          ack1 => if_stmt_615_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_822_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond22_821;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_822_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_822_branch_req_0,
          ack0 => if_stmt_822_branch_ack_0,
          ack1 => if_stmt_822_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_837_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264448_836;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_837_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_837_branch_req_0,
          ack0 => if_stmt_837_branch_ack_0,
          ack1 => if_stmt_837_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_912_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_911;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_912_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_912_branch_req_0,
          ack0 => if_stmt_912_branch_ack_0,
          ack1 => if_stmt_912_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1001_inst
    process(input_dim2_966, nao2_997) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2_966, nao2_997, tmp_var);
      nao3_1002 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1067_inst
    process(input_dim2_966) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2_966, konst_1066_wire_constant, tmp_var);
      nid2_true_1068 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1072_inst
    process(input_dim1_962) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1_962, konst_1071_wire_constant, tmp_var);
      nid2_false_1073 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1077_inst
    process(add_dest_dim1_974, stride_226) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_dest_dim1_974, stride_226, tmp_var);
      nid2_false1_1078 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1082_inst
    process(input_dim0_958) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0_958, konst_1081_wire_constant, tmp_var);
      nid1_true_1083 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1087_inst
    process(add_dest_dim0_970, stride_226) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_dest_dim0_970, stride_226, tmp_var);
      nid1_true1_1088 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_940_inst
    process(padding_251) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(padding_251, konst_939_wire_constant, tmp_var);
      pad_941 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_991_inst
    process(nao_987, add_dest_dim1_974) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nao_987, add_dest_dim1_974, tmp_var);
      nao1_992 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1110_inst
    process(add_src_978) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_src_978, konst_1109_wire_constant, tmp_var);
      next_add_src_1111 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1316_inst
    process(tmp464_1305) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp464_1305, type_cast_1315_wire_constant, tmp_var);
      tmp464x_xop_1317 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_431_inst
    process(tmp495_420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp495_420, type_cast_430_wire_constant, tmp_var);
      tmp495x_xop_432 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_638_inst
    process(tmp482_627) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp482_627, type_cast_637_wire_constant, tmp_var);
      tmp482x_xop_639 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_860_inst
    process(tmp476_849) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp476_849, type_cast_859_wire_constant, tmp_var);
      tmp476x_xop_861 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1326_inst
    process(iNsTr_111_1321) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_111_1321, type_cast_1325_wire_constant, tmp_var);
      xx_xop_1327 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1458_inst
    process(indvar_1337) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1337, type_cast_1457_wire_constant, tmp_var);
      indvarx_xnext_1459 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_441_inst
    process(iNsTr_19_436) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_19_436, type_cast_440_wire_constant, tmp_var);
      xx_xop503_442 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_608_inst
    process(indvar489_452) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar489_452, type_cast_607_wire_constant, tmp_var);
      indvarx_xnext490_609 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_648_inst
    process(iNsTr_32_643) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_32_643, type_cast_647_wire_constant, tmp_var);
      xx_xop502_649 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_815_inst
    process(indvar476_659) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar476_659, type_cast_814_wire_constant, tmp_var);
      indvarx_xnext477_816 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_870_inst
    process(iNsTr_52_865) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_52_865, type_cast_869_wire_constant, tmp_var);
      xx_xop513_871 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_905_inst
    process(indvar469_881) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar469_881, type_cast_904_wire_constant, tmp_var);
      indvarx_xnext470_906 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1062_inst
    process(NOT_u1_u1_1060_wire, cmp_dim1_1057) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1060_wire, cmp_dim1_1057, tmp_var);
      cmp_dim0_1063 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1056_inst
    process(input_dim1_962, SUB_u16_u16_1046_1046_delayed_1_0_1052) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim1_962, SUB_u16_u16_1046_1046_delayed_1_0_1052, tmp_var);
      cmp_dim1_1057 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1463_inst
    process(indvarx_xnext_1459, tmp468_1334) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1459, tmp468_1334, tmp_var);
      exitcond1_1464 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_613_inst
    process(indvarx_xnext490_609, tmp500_449) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext490_609, tmp500_449, tmp_var);
      exitcond2_614 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_820_inst
    process(indvarx_xnext477_816, tmp487_656) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext477_816, tmp487_656, tmp_var);
      exitcond22_821 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_910_inst
    process(indvarx_xnext470_906, tmp481_878) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext470_906, tmp481_878, tmp_var);
      exitcond_911 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1006_inst
    process(nao3_1002) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nao3_1002, konst_1005_wire_constant, tmp_var);
      add_out_1007 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1304_inst
    process(output_size_386) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(output_size_386, type_cast_1303_wire_constant, tmp_var);
      tmp464_1305 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_419_inst
    process(input_size_345) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(input_size_345, type_cast_418_wire_constant, tmp_var);
      tmp495_420 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_626_inst
    process(kernel_size_368) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(kernel_size_368, type_cast_625_wire_constant, tmp_var);
      tmp482_627 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_848_inst
    process(output_size_386) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(output_size_386, type_cast_847_wire_constant, tmp_var);
      tmp476_849 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1196_inst
    process(sub_1186) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1186, type_cast_1195_wire_constant, tmp_var);
      shr308_1197 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1206_inst
    process(sub_1186) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1186, type_cast_1205_wire_constant, tmp_var);
      shr314_1207 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1216_inst
    process(sub_1186) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1186, type_cast_1215_wire_constant, tmp_var);
      shr320_1217 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1226_inst
    process(sub_1186) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1186, type_cast_1225_wire_constant, tmp_var);
      shr326_1227 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1236_inst
    process(sub_1186) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1186, type_cast_1235_wire_constant, tmp_var);
      shr332_1237 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1246_inst
    process(sub_1186) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1186, type_cast_1245_wire_constant, tmp_var);
      shr338_1247 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1256_inst
    process(sub_1186) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1186, type_cast_1255_wire_constant, tmp_var);
      shr344_1257 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1364_inst
    process(tmp377_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_1355, type_cast_1363_wire_constant, tmp_var);
      shr384_1365 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1374_inst
    process(tmp377_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_1355, type_cast_1373_wire_constant, tmp_var);
      shr390_1375 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1384_inst
    process(tmp377_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_1355, type_cast_1383_wire_constant, tmp_var);
      shr396_1385 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1394_inst
    process(tmp377_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_1355, type_cast_1393_wire_constant, tmp_var);
      shr402_1395 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1404_inst
    process(tmp377_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_1355, type_cast_1403_wire_constant, tmp_var);
      shr408_1405 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1414_inst
    process(tmp377_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_1355, type_cast_1413_wire_constant, tmp_var);
      shr414_1415 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1424_inst
    process(tmp377_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp377_1355, type_cast_1423_wire_constant, tmp_var);
      shr420_1425 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1092_inst
    process(stride_226, inp_d1_76) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(stride_226, inp_d1_76, tmp_var);
      nid1_true2_1093 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_335_inst
    process(inp_d0_51, inp_d1_76) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(inp_d0_51, inp_d1_76, tmp_var);
      input_int_336 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_349_inst
    process(ker_d0_126, ker_d1_151) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ker_d0_126, ker_d1_151, tmp_var);
      ker_int1_350 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_354_inst
    process(ker_d2_176, ker_d3_201) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ker_d2_176, ker_d3_201, tmp_var);
      ker_int2_355 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_376_inst
    process(out_d0_276, out_d1_301) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_d0_276, out_d1_301, tmp_var);
      out_int_377 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_986_inst
    process(out_d1_301, add_dest_dim0_970) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_d1_301, add_dest_dim0_970, tmp_var);
      nao_987 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_996_inst
    process(out_d2_326, nao1_992) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_d2_326, nao1_992, tmp_var);
      nao2_997 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_344_inst
    process(input_int1_340, inp_d232_331) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_int1_340, inp_d232_331, tmp_var);
      input_size_345 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_367_inst
    process(ker_int3_359, ker_int4_363) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(ker_int3_359, ker_int4_363, tmp_var);
      kernel_size_368 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_385_inst
    process(out_int1_381, out_d232_372) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(out_int1_381, out_d232_372, tmp_var);
      output_size_386 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1060_inst
    process(cmp_dim2_1047) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_1047, tmp_var);
      NOT_u1_u1_1060_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1114_inst
    process(cmp_dim2_1047) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_1047, tmp_var);
      NOT_u1_u1_1114_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1136_inst
    process(cmp_dim2_1047) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim2_1047, tmp_var);
      NOT_u1_u1_1136_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1163_inst
    process(cmp_dim0_1063) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_dim0_1063, tmp_var);
      NOT_u1_u1_1163_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_100_inst
    process(shl18_89, conv20_96) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_89, conv20_96, tmp_var);
      inp_d2_101 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_125_inst
    process(shl27_114, conv29_121) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_114, conv29_121, tmp_var);
      ker_d0_126 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_150_inst
    process(shl36_139, conv38_146) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_139, conv38_146, tmp_var);
      ker_d1_151 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_175_inst
    process(shl45_164, conv47_171) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_164, conv47_171, tmp_var);
      ker_d2_176 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_200_inst
    process(shl54_189, conv56_196) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_189, conv56_196, tmp_var);
      ker_d3_201 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_225_inst
    process(shl96_214, conv98_221) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_214, conv98_221, tmp_var);
      stride_226 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_250_inst
    process(shl105_239, conv107_246) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_239, conv107_246, tmp_var);
      padding_251 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_275_inst
    process(shl114_264, conv116_271) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_264, conv116_271, tmp_var);
      out_d0_276 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_300_inst
    process(shl123_289, conv1125_296) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_289, conv1125_296, tmp_var);
      out_d1_301 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_325_inst
    process(shl132_314, conv134_321) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_314, conv134_321, tmp_var);
      out_d2_326 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_50_inst
    process(shl_39, conv3_46) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_39, conv3_46, tmp_var);
      inp_d0_51 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_75_inst
    process(shl9_64, conv11_71) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_64, conv11_71, tmp_var);
      inp_d1_76 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1164_inst
    process(dim0_end_1159, NOT_u1_u1_1163_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(dim0_end_1159, NOT_u1_u1_1163_wire, tmp_var);
      continue_flag_1165 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_490_inst
    process(shl127_479, conv130_486) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl127_479, conv130_486, tmp_var);
      add131_491 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_508_inst
    process(shl133_497, conv136_504) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl133_497, conv136_504, tmp_var);
      add137_509 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_526_inst
    process(shl139_515, conv142_522) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl139_515, conv142_522, tmp_var);
      add143_527 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_544_inst
    process(shl145_533, conv148_540) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl145_533, conv148_540, tmp_var);
      add149_545 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_562_inst
    process(shl151_551, conv154_558) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl151_551, conv154_558, tmp_var);
      add155_563 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_580_inst
    process(shl157_569, conv160_576) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl157_569, conv160_576, tmp_var);
      add161_581 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_598_inst
    process(shl163_587, conv166_594) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl163_587, conv166_594, tmp_var);
      add167_599 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_697_inst
    process(shl183_686, conv186_693) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl183_686, conv186_693, tmp_var);
      add187_698 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_715_inst
    process(shl189_704, conv192_711) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl189_704, conv192_711, tmp_var);
      add193_716 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_733_inst
    process(shl195_722, conv198_729) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl195_722, conv198_729, tmp_var);
      add199_734 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_751_inst
    process(shl201_740, conv204_747) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl201_740, conv204_747, tmp_var);
      add205_752 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_769_inst
    process(shl207_758, conv210_765) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl207_758, conv210_765, tmp_var);
      add211_770 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_787_inst
    process(shl213_776, conv216_783) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl213_776, conv216_783, tmp_var);
      add217_788 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_805_inst
    process(shl219_794, conv222_801) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl219_794, conv222_801, tmp_var);
      add223_806 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_113_inst
    process(conv26_108) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_108, type_cast_112_wire_constant, tmp_var);
      shl27_114 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_138_inst
    process(conv35_133) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_133, type_cast_137_wire_constant, tmp_var);
      shl36_139 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_163_inst
    process(conv44_158) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_158, type_cast_162_wire_constant, tmp_var);
      shl45_164 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_188_inst
    process(conv53_183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_183, type_cast_187_wire_constant, tmp_var);
      shl54_189 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_213_inst
    process(conv95_208) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_208, type_cast_212_wire_constant, tmp_var);
      shl96_214 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_238_inst
    process(conv104_233) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_233, type_cast_237_wire_constant, tmp_var);
      shl105_239 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_263_inst
    process(conv113_258) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_258, type_cast_262_wire_constant, tmp_var);
      shl114_264 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_288_inst
    process(conv122_283) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_283, type_cast_287_wire_constant, tmp_var);
      shl123_289 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_313_inst
    process(conv131_308) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_308, type_cast_312_wire_constant, tmp_var);
      shl132_314 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_38_inst
    process(conv1_33) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_33, type_cast_37_wire_constant, tmp_var);
      shl_39 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_63_inst
    process(conv8_58) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_58, type_cast_62_wire_constant, tmp_var);
      shl9_64 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_88_inst
    process(conv17_83) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_83, type_cast_87_wire_constant, tmp_var);
      shl18_89 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_478_inst
    process(conv125_473) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv125_473, type_cast_477_wire_constant, tmp_var);
      shl127_479 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_496_inst
    process(add131_491) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add131_491, type_cast_495_wire_constant, tmp_var);
      shl133_497 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_514_inst
    process(add137_509) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add137_509, type_cast_513_wire_constant, tmp_var);
      shl139_515 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_532_inst
    process(add143_527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add143_527, type_cast_531_wire_constant, tmp_var);
      shl145_533 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_550_inst
    process(add149_545) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add149_545, type_cast_549_wire_constant, tmp_var);
      shl151_551 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_568_inst
    process(add155_563) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add155_563, type_cast_567_wire_constant, tmp_var);
      shl157_569 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_586_inst
    process(add161_581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add161_581, type_cast_585_wire_constant, tmp_var);
      shl163_587 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_685_inst
    process(conv181_680) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv181_680, type_cast_684_wire_constant, tmp_var);
      shl183_686 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_703_inst
    process(add187_698) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add187_698, type_cast_702_wire_constant, tmp_var);
      shl189_704 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_721_inst
    process(add193_716) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add193_716, type_cast_720_wire_constant, tmp_var);
      shl195_722 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_739_inst
    process(add199_734) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add199_734, type_cast_738_wire_constant, tmp_var);
      shl201_740 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_757_inst
    process(add205_752) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add205_752, type_cast_756_wire_constant, tmp_var);
      shl207_758 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_775_inst
    process(add211_770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add211_770, type_cast_774_wire_constant, tmp_var);
      shl213_776 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_793_inst
    process(add217_788) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add217_788, type_cast_792_wire_constant, tmp_var);
      shl219_794 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1038_inst
    process(inp_d2_101) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(inp_d2_101, konst_1037_wire_constant, tmp_var);
      dim2_limit_1039 <= tmp_var; --
    end process;
    -- shared split operator group (114) : SUB_u16_u16_1051_inst 
    ApIntSub_group_114: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= inp_d1_76;
      SUB_u16_u16_1046_1046_delayed_1_0_1052 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_1051_inst_req_0;
      SUB_u16_u16_1051_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_1051_inst_req_1;
      SUB_u16_u16_1051_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_114_gI: SplitGuardInterface generic map(name => "ApIntSub_group_114_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_114",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 114
    -- binary operator SUB_u16_u16_1097_inst
    process(nid1_true2_1093, stride_226) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(nid1_true2_1093, stride_226, tmp_var);
      nid1_true3_1098 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1105_inst
    process(add_dest_dim1_974, nid1_true3_1092_delayed_1_0_1101) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add_dest_dim1_974, nid1_true3_1092_delayed_1_0_1101, tmp_var);
      nid1_true4_1106 <= tmp_var; --
    end process;
    -- shared split operator group (117) : SUB_u16_u16_1153_inst 
    ApIntSub_group_117: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= inp_d0_51;
      SUB_u16_u16_1142_1142_delayed_1_0_1154 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_1153_inst_req_0;
      SUB_u16_u16_1153_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_1153_inst_req_1;
      SUB_u16_u16_1153_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_117_gI: SplitGuardInterface generic map(name => "ApIntSub_group_117_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- binary operator SUB_u16_u16_945_inst
    process(ker_d1_151, pad_941) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(ker_d1_151, pad_941, tmp_var);
      add_dest_dim0_init_946 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_950_inst
    process(ker_d2_176, pad_941) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(ker_d2_176, pad_941, tmp_var);
      add_dest_dim1_init_951 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1185_inst
    process(conv298_1181, conv276_1176) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv298_1181, conv276_1176, tmp_var);
      sub_1186 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1291_inst
    process(output_size_386) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(output_size_386, type_cast_1290_wire_constant, tmp_var);
      cmp264449_1292 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1310_inst
    process(tmp464_1305) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp464_1305, type_cast_1309_wire_constant, tmp_var);
      tmp465_1311 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_391_inst
    process(input_size_345) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(input_size_345, type_cast_390_wire_constant, tmp_var);
      cmp467_392 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_406_inst
    process(kernel_size_368) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(kernel_size_368, type_cast_405_wire_constant, tmp_var);
      cmp175463_407 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_425_inst
    process(tmp495_420) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp495_420, type_cast_424_wire_constant, tmp_var);
      tmp496_426 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_632_inst
    process(tmp482_627) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp482_627, type_cast_631_wire_constant, tmp_var);
      tmp483_633 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_835_inst
    process(output_size_386) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(output_size_386, type_cast_834_wire_constant, tmp_var);
      cmp264448_836 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_854_inst
    process(tmp476_849) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp476_849, type_cast_853_wire_constant, tmp_var);
      tmp477_855 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_1046_inst
    process(input_dim2_966, dim2_limit_1039_delayed_1_0_1042) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(input_dim2_966, dim2_limit_1039_delayed_1_0_1042, tmp_var);
      cmp_dim2_1047 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_1158_inst
    process(input_dim0_958, SUB_u16_u16_1142_1142_delayed_1_0_1154) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(input_dim0_958, SUB_u16_u16_1142_1142_delayed_1_0_1154, tmp_var);
      dim0_end_1159 <= tmp_var; --
    end process;
    -- shared split operator group (131) : array_obj_ref_1013_index_offset 
    ApIntAdd_group_131: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_1012_scaled;
      array_obj_ref_1013_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1013_index_offset_req_0;
      array_obj_ref_1013_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1013_index_offset_req_1;
      array_obj_ref_1013_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_131_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_131_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_131",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 131
    -- shared split operator group (132) : array_obj_ref_1025_index_offset 
    ApIntAdd_group_132: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_1024_scaled;
      array_obj_ref_1025_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1025_index_offset_req_0;
      array_obj_ref_1025_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1025_index_offset_req_1;
      array_obj_ref_1025_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_132_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_132_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_132",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 132
    -- shared split operator group (133) : array_obj_ref_1349_index_offset 
    ApIntAdd_group_133: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1348_scaled;
      array_obj_ref_1349_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1349_index_offset_req_0;
      array_obj_ref_1349_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1349_index_offset_req_1;
      array_obj_ref_1349_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_133_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_133_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_133",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 133
    -- shared split operator group (134) : array_obj_ref_464_index_offset 
    ApIntAdd_group_134: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar489_463_scaled;
      array_obj_ref_464_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_464_index_offset_req_0;
      array_obj_ref_464_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_464_index_offset_req_1;
      array_obj_ref_464_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_134_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_134_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_134",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 134
    -- shared split operator group (135) : array_obj_ref_671_index_offset 
    ApIntAdd_group_135: Block -- 
      signal data_in: std_logic_vector(9 downto 0);
      signal data_out: std_logic_vector(9 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar476_670_scaled;
      array_obj_ref_671_final_offset <= data_out(9 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_671_index_offset_req_0;
      array_obj_ref_671_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_671_index_offset_req_1;
      array_obj_ref_671_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_135_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_135_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_135",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 10,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 10,
          constant_operand => "0000000000",
          constant_width => 10,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 135
    -- shared split operator group (136) : array_obj_ref_893_index_offset 
    ApIntAdd_group_136: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar469_892_scaled;
      array_obj_ref_893_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_893_index_offset_req_0;
      array_obj_ref_893_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_893_index_offset_req_1;
      array_obj_ref_893_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_136_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_136_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_136",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 136
    -- unary operator type_cast_1174_inst
    process(call233_923) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call233_923, tmp_var);
      type_cast_1174_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1179_inst
    process(call297_1170) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call297_1170, tmp_var);
      type_cast_1179_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1018_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1018_load_0_req_0;
      ptr_deref_1018_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1018_load_0_req_1;
      ptr_deref_1018_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1018_word_address_0;
      ptr_deref_1018_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1354_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1354_load_0_req_0;
      ptr_deref_1354_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1354_load_0_req_1;
      ptr_deref_1354_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1354_word_address_0;
      ptr_deref_1354_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : ptr_deref_1032_store_0 ptr_deref_897_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1032_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_897_store_0_req_0;
      ptr_deref_1032_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_897_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1032_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_897_store_0_req_1;
      ptr_deref_1032_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_897_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1032_word_address_0 & ptr_deref_897_word_address_0;
      data_in <= ptr_deref_1032_data_0 & ptr_deref_897_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_601_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_601_store_0_req_0;
      ptr_deref_601_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_601_store_0_req_1;
      ptr_deref_601_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_601_word_address_0;
      data_in <= ptr_deref_601_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_808_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(9 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_808_store_0_req_0;
      ptr_deref_808_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_808_store_0_req_1;
      ptr_deref_808_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_808_word_address_0;
      data_in <= ptr_deref_808_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 10,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(9 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_778_inst RPIPE_ConvTranspose_input_pipe_742_inst RPIPE_ConvTranspose_input_pipe_675_inst RPIPE_ConvTranspose_input_pipe_688_inst RPIPE_ConvTranspose_input_pipe_724_inst RPIPE_ConvTranspose_input_pipe_796_inst RPIPE_ConvTranspose_input_pipe_706_inst RPIPE_ConvTranspose_input_pipe_760_inst RPIPE_ConvTranspose_input_pipe_166_inst RPIPE_ConvTranspose_input_pipe_153_inst RPIPE_ConvTranspose_input_pipe_216_inst RPIPE_ConvTranspose_input_pipe_27_inst RPIPE_ConvTranspose_input_pipe_116_inst RPIPE_ConvTranspose_input_pipe_228_inst RPIPE_ConvTranspose_input_pipe_103_inst RPIPE_ConvTranspose_input_pipe_241_inst RPIPE_ConvTranspose_input_pipe_91_inst RPIPE_ConvTranspose_input_pipe_203_inst RPIPE_ConvTranspose_input_pipe_178_inst RPIPE_ConvTranspose_input_pipe_78_inst RPIPE_ConvTranspose_input_pipe_141_inst RPIPE_ConvTranspose_input_pipe_128_inst RPIPE_ConvTranspose_input_pipe_66_inst RPIPE_ConvTranspose_input_pipe_191_inst RPIPE_ConvTranspose_input_pipe_53_inst RPIPE_ConvTranspose_input_pipe_41_inst RPIPE_ConvTranspose_input_pipe_253_inst RPIPE_ConvTranspose_input_pipe_266_inst RPIPE_ConvTranspose_input_pipe_278_inst RPIPE_ConvTranspose_input_pipe_291_inst RPIPE_ConvTranspose_input_pipe_303_inst RPIPE_ConvTranspose_input_pipe_316_inst RPIPE_ConvTranspose_input_pipe_468_inst RPIPE_ConvTranspose_input_pipe_481_inst RPIPE_ConvTranspose_input_pipe_499_inst RPIPE_ConvTranspose_input_pipe_517_inst RPIPE_ConvTranspose_input_pipe_535_inst RPIPE_ConvTranspose_input_pipe_553_inst RPIPE_ConvTranspose_input_pipe_571_inst RPIPE_ConvTranspose_input_pipe_589_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_778_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_742_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_675_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_688_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_724_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_796_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_706_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_760_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_166_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_153_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_216_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_27_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_116_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_228_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_103_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_241_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_91_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_203_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_178_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_78_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_141_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_66_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_191_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_41_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_253_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_266_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_278_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_291_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_303_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_468_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_481_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_499_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_517_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_535_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_553_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_571_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_589_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_778_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_742_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_675_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_688_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_724_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_796_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_706_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_760_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_166_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_153_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_216_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_27_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_116_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_228_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_103_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_241_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_91_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_203_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_178_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_78_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_141_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_66_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_191_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_41_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_253_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_266_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_278_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_291_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_303_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_468_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_481_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_499_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_517_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_535_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_553_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_571_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_589_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_778_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_742_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_675_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_688_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_724_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_796_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_706_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_760_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_166_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_153_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_216_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_27_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_116_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_228_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_103_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_241_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_91_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_203_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_178_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_78_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_141_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_66_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_191_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_41_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_253_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_266_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_278_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_291_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_303_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_468_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_481_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_499_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_517_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_535_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_553_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_571_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_589_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_778_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_742_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_675_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_688_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_724_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_796_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_706_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_760_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_166_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_153_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_216_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_27_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_116_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_228_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_103_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_241_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_91_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_203_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_178_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_78_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_141_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_66_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_191_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_41_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_253_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_266_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_278_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_291_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_303_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_468_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_481_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_499_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_517_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_535_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_553_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_571_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_589_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call214_779 <= data_out(319 downto 312);
      call202_743 <= data_out(311 downto 304);
      call180_676 <= data_out(303 downto 296);
      call184_689 <= data_out(295 downto 288);
      call196_725 <= data_out(287 downto 280);
      call220_797 <= data_out(279 downto 272);
      call190_707 <= data_out(271 downto 264);
      call208_761 <= data_out(263 downto 256);
      call46_167 <= data_out(255 downto 248);
      call41_154 <= data_out(247 downto 240);
      call97_217 <= data_out(239 downto 232);
      call_28 <= data_out(231 downto 224);
      call28_117 <= data_out(223 downto 216);
      call101_229 <= data_out(215 downto 208);
      call23_104 <= data_out(207 downto 200);
      call106_242 <= data_out(199 downto 192);
      call19_92 <= data_out(191 downto 184);
      call92_204 <= data_out(183 downto 176);
      call50_179 <= data_out(175 downto 168);
      call14_79 <= data_out(167 downto 160);
      call37_142 <= data_out(159 downto 152);
      call32_129 <= data_out(151 downto 144);
      call10_67 <= data_out(143 downto 136);
      call55_192 <= data_out(135 downto 128);
      call5_54 <= data_out(127 downto 120);
      call2_42 <= data_out(119 downto 112);
      call110_254 <= data_out(111 downto 104);
      call115_267 <= data_out(103 downto 96);
      call119_279 <= data_out(95 downto 88);
      call1124_292 <= data_out(87 downto 80);
      call1128_304 <= data_out(79 downto 72);
      call133_317 <= data_out(71 downto 64);
      call124_469 <= data_out(63 downto 56);
      call128_482 <= data_out(55 downto 48);
      call134_500 <= data_out(47 downto 40);
      call140_518 <= data_out(39 downto 32);
      call146_536 <= data_out(31 downto 24);
      call152_554 <= data_out(23 downto 16);
      call158_572 <= data_out(15 downto 8);
      call164_590 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_1274_inst WPIPE_ConvTranspose_output_pipe_1277_inst WPIPE_ConvTranspose_output_pipe_1262_inst WPIPE_ConvTranspose_output_pipe_1280_inst WPIPE_ConvTranspose_output_pipe_1268_inst WPIPE_ConvTranspose_output_pipe_1283_inst WPIPE_ConvTranspose_output_pipe_1265_inst WPIPE_ConvTranspose_output_pipe_1271_inst WPIPE_ConvTranspose_output_pipe_1430_inst WPIPE_ConvTranspose_output_pipe_1433_inst WPIPE_ConvTranspose_output_pipe_1436_inst WPIPE_ConvTranspose_output_pipe_1439_inst WPIPE_ConvTranspose_output_pipe_1442_inst WPIPE_ConvTranspose_output_pipe_1445_inst WPIPE_ConvTranspose_output_pipe_1448_inst WPIPE_ConvTranspose_output_pipe_1451_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1274_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1277_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1262_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1280_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1268_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1283_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1265_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1271_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1430_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1433_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1436_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1439_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1442_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1445_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1448_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1451_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1274_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1277_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1262_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1280_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1268_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1283_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1265_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1271_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1430_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1433_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1436_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1439_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1442_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1445_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1274_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1277_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1262_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1280_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1268_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1283_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1265_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1271_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1430_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1433_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1436_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1439_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1442_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1445_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1448_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1451_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1274_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1277_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1262_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1280_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1268_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1283_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1265_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1271_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1430_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1433_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1436_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1439_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1442_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1445_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv323_1221 & conv317_1211 & conv347_1261 & conv311_1201 & conv335_1241 & conv305_1191 & conv341_1251 & conv329_1231 & conv423_1429 & conv417_1419 & conv411_1409 & conv405_1399 & conv399_1389 & conv393_1379 & conv387_1369 & conv381_1359;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_923_call call_stmt_1170_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_923_call_req_0;
      reqL_unguarded(0) <= call_stmt_1170_call_req_0;
      call_stmt_923_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1170_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_923_call_req_1;
      reqR_unguarded(0) <= call_stmt_1170_call_req_1;
      call_stmt_923_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1170_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call233_923 <= data_out(127 downto 64);
      call297_1170 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end ct_core_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_16_inst_req_0 : boolean;
  signal WPIPE_timer_req_16_inst_ack_0 : boolean;
  signal WPIPE_timer_req_16_inst_req_1 : boolean;
  signal WPIPE_timer_req_16_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_21_inst_req_0 : boolean;
  signal RPIPE_timer_resp_21_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_21_inst_req_1 : boolean;
  signal RPIPE_timer_resp_21_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_19_to_assign_stmt_22/$entry
      -- CP-element group 0: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_sample_start_
      -- CP-element group 0: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_Sample/req
      -- CP-element group 0: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_sample_start_
      -- CP-element group 0: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_Sample/rr
      -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_21_inst_req_0); -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_16_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_sample_completed_
      -- CP-element group 1: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_update_start_
      -- CP-element group 1: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_Sample/ack
      -- CP-element group 1: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_Update/$entry
      -- CP-element group 1: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_16_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_16_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_update_completed_
      -- CP-element group 2: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_Update/$exit
      -- CP-element group 2: 	 assign_stmt_19_to_assign_stmt_22/WPIPE_timer_req_16_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_16_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_update_start_
      -- CP-element group 3: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_sample_completed_
      -- CP-element group 3: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_Sample/ra
      -- CP-element group 3: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_Update/$entry
      -- CP-element group 3: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_21_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_21_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_update_completed_
      -- CP-element group 4: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_Update/$exit
      -- CP-element group 4: 	 assign_stmt_19_to_assign_stmt_22/RPIPE_timer_resp_21_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_21_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_19_to_assign_stmt_22/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(4) & timer_CP_0_elements(2);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_18_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_18_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_21_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_21_inst_req_0;
      RPIPE_timer_resp_21_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_21_inst_req_1;
      RPIPE_timer_resp_21_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_16_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_16_inst_req_0;
      WPIPE_timer_req_16_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_16_inst_req_1;
      WPIPE_timer_req_16_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_18_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_3369_start: Boolean;
  signal timerDaemon_CP_3369_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_timer_req_1492_inst_req_0 : boolean;
  signal RPIPE_timer_req_1492_inst_req_1 : boolean;
  signal RPIPE_timer_req_1492_inst_ack_0 : boolean;
  signal RPIPE_timer_req_1492_inst_ack_1 : boolean;
  signal nCOUNTER_1498_1489_buf_ack_1 : boolean;
  signal do_while_stmt_1483_branch_ack_0 : boolean;
  signal do_while_stmt_1483_branch_ack_1 : boolean;
  signal nCOUNTER_1498_1489_buf_req_1 : boolean;
  signal phi_stmt_1485_req_0 : boolean;
  signal WPIPE_timer_resp_1500_inst_req_0 : boolean;
  signal WPIPE_timer_resp_1500_inst_ack_0 : boolean;
  signal nCOUNTER_1498_1489_buf_ack_0 : boolean;
  signal phi_stmt_1485_req_1 : boolean;
  signal nCOUNTER_1498_1489_buf_req_0 : boolean;
  signal phi_stmt_1485_ack_0 : boolean;
  signal WPIPE_timer_resp_1500_inst_req_1 : boolean;
  signal WPIPE_timer_resp_1500_inst_ack_1 : boolean;
  signal do_while_stmt_1483_branch_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_3369_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3369_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_3369_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3369_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_3369: Block -- control-path 
    signal timerDaemon_CP_3369_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_3369_elements(0) <= timerDaemon_CP_3369_start;
    timerDaemon_CP_3369_symbol <= timerDaemon_CP_3369_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1482/branch_block_stmt_1482__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1482/do_while_stmt_1483__entry__
      -- CP-element group 0: 	 branch_block_stmt_1482/$entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1482/do_while_stmt_1483__exit__
      -- CP-element group 1: 	 branch_block_stmt_1482/branch_block_stmt_1482__exit__
      -- CP-element group 1: 	 branch_block_stmt_1482/$exit
      -- CP-element group 1: 	 $exit
      -- 
    timerDaemon_CP_3369_elements(1) <= timerDaemon_CP_3369_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1482/do_while_stmt_1483/$entry
      -- CP-element group 2: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483__entry__
      -- 
    timerDaemon_CP_3369_elements(2) <= timerDaemon_CP_3369_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483__exit__
      -- 
    -- Element group timerDaemon_CP_3369_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1482/do_while_stmt_1483/loop_back
      -- 
    -- Element group timerDaemon_CP_3369_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1482/do_while_stmt_1483/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1482/do_while_stmt_1483/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1482/do_while_stmt_1483/loop_taken/$entry
      -- 
    timerDaemon_CP_3369_elements(5) <= timerDaemon_CP_3369_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1482/do_while_stmt_1483/loop_body_done
      -- 
    timerDaemon_CP_3369_elements(6) <= timerDaemon_CP_3369_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_3369_elements(7) <= timerDaemon_CP_3369_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_3369_elements(8) <= timerDaemon_CP_3369_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1490_sample_start_
      -- 
    -- Element group timerDaemon_CP_3369_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	40 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/condition_evaluated
      -- 
    condition_evaluated_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3369_elements(10), ack => do_while_stmt_1483_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(14) & timerDaemon_CP_3369_elements(40);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(9) & timerDaemon_CP_3369_elements(15) & timerDaemon_CP_3369_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1490_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(17) & timerDaemon_CP_3369_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(16) & timerDaemon_CP_3369_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(18) & timerDaemon_CP_3369_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(9) & timerDaemon_CP_3369_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(9) & timerDaemon_CP_3369_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_3369_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_update_completed_
      -- 
    -- Element group timerDaemon_CP_3369_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_loopback_trigger
      -- 
    timerDaemon_CP_3369_elements(19) <= timerDaemon_CP_3369_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_loopback_sample_req_ps
      -- 
    phi_stmt_1485_loopback_sample_req_3408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1485_loopback_sample_req_3408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3369_elements(20), ack => phi_stmt_1485_req_1); -- 
    -- Element group timerDaemon_CP_3369_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_entry_trigger
      -- 
    timerDaemon_CP_3369_elements(21) <= timerDaemon_CP_3369_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_entry_sample_req
      -- 
    phi_stmt_1485_entry_sample_req_3411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1485_entry_sample_req_3411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3369_elements(22), ack => phi_stmt_1485_req_0); -- 
    -- Element group timerDaemon_CP_3369_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1485_phi_mux_ack_ps
      -- 
    phi_stmt_1485_phi_mux_ack_3414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1485_ack_0, ack => timerDaemon_CP_3369_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/type_cast_1488_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/type_cast_1488_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/type_cast_1488_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/type_cast_1488_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_3369_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/type_cast_1488_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/type_cast_1488_update_start__ps
      -- 
    -- Element group timerDaemon_CP_3369_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/type_cast_1488_update_completed__ps
      -- 
    timerDaemon_CP_3369_elements(26) <= timerDaemon_CP_3369_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/type_cast_1488_update_completed_
      -- 
    -- Element group timerDaemon_CP_3369_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_3369_elements(25), ack => timerDaemon_CP_3369_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_sample_start_
      -- 
    req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3369_elements(28), ack => nCOUNTER_1498_1489_buf_req_0); -- 
    -- Element group timerDaemon_CP_3369_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_Update/req
      -- CP-element group 29: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_update_start_
      -- 
    req_3440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3369_elements(29), ack => nCOUNTER_1498_1489_buf_req_1); -- 
    -- Element group timerDaemon_CP_3369_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_Sample/$exit
      -- 
    ack_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1498_1489_buf_ack_0, ack => timerDaemon_CP_3369_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/R_nCOUNTER_1489_update_completed_
      -- 
    ack_3441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1498_1489_buf_ack_1, ack => timerDaemon_CP_3369_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1490_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(9) & timerDaemon_CP_3369_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_sample_start_
      -- 
    rr_3454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3369_elements(33), ack => RPIPE_timer_req_1492_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(11) & timerDaemon_CP_3369_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_Update/$entry
      -- 
    cr_3459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3369_elements(34), ack => RPIPE_timer_req_1492_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(13) & timerDaemon_CP_3369_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_Sample/$exit
      -- 
    ra_3455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1492_inst_ack_0, ack => timerDaemon_CP_3369_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/phi_stmt_1490_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/RPIPE_timer_req_1492_update_completed_
      -- 
    ca_3460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1492_inst_ack_1, ack => timerDaemon_CP_3369_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_Sample/req
      -- 
    req_3468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3369_elements(37), ack => WPIPE_timer_resp_1500_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(18) & timerDaemon_CP_3369_elements(36) & timerDaemon_CP_3369_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_Update/req
      -- 
    ack_3469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1500_inst_ack_0, ack => timerDaemon_CP_3369_elements(38)); -- 
    req_3473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3369_elements(38), ack => WPIPE_timer_resp_1500_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/WPIPE_timer_resp_1500_Update/ack
      -- 
    ack_3474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1500_inst_ack_1, ack => timerDaemon_CP_3369_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_3369_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_3369_elements(9), ack => timerDaemon_CP_3369_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1482/do_while_stmt_1483/do_while_stmt_1483_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3369_elements(12) & timerDaemon_CP_3369_elements(39);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3369_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1482/do_while_stmt_1483/loop_exit/ack
      -- CP-element group 42: 	 branch_block_stmt_1482/do_while_stmt_1483/loop_exit/$exit
      -- 
    ack_3479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1483_branch_ack_0, ack => timerDaemon_CP_3369_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1482/do_while_stmt_1483/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_1482/do_while_stmt_1483/loop_taken/ack
      -- 
    ack_3483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1483_branch_ack_1, ack => timerDaemon_CP_3369_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1482/do_while_stmt_1483/$exit
      -- 
    timerDaemon_CP_3369_elements(44) <= timerDaemon_CP_3369_elements(3);
    timerDaemon_do_while_stmt_1483_terminator_3484: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1483_terminator_3484", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_3369_elements(6),loop_continue => timerDaemon_CP_3369_elements(43),loop_terminate => timerDaemon_CP_3369_elements(42),loop_back => timerDaemon_CP_3369_elements(4),loop_exit => timerDaemon_CP_3369_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1485_phi_seq_3442_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_3369_elements(21);
      timerDaemon_CP_3369_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_3369_elements(24);
      timerDaemon_CP_3369_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_3369_elements(26);
      timerDaemon_CP_3369_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_3369_elements(19);
      timerDaemon_CP_3369_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_3369_elements(30);
      timerDaemon_CP_3369_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_3369_elements(31);
      timerDaemon_CP_3369_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1485_phi_seq_3442 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1485_phi_seq_3442") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_3369_elements(11), 
          phi_sample_ack => timerDaemon_CP_3369_elements(17), 
          phi_update_req => timerDaemon_CP_3369_elements(13), 
          phi_update_ack => timerDaemon_CP_3369_elements(18), 
          phi_mux_ack => timerDaemon_CP_3369_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3394_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_3369_elements(7);
        preds(1)  <= timerDaemon_CP_3369_elements(8);
        entry_tmerge_3394 : transition_merge -- 
          generic map(name => " entry_tmerge_3394")
          port map (preds => preds, symbol_out => timerDaemon_CP_3369_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_1485 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_1492_wire : std_logic_vector(0 downto 0);
    signal konst_1496_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1504_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_1498 : std_logic_vector(63 downto 0);
    signal nCOUNTER_1498_1489_buffered : std_logic_vector(63 downto 0);
    signal req_1490 : std_logic_vector(0 downto 0);
    signal type_cast_1488_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1496_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1504_wire_constant <= "1";
    type_cast_1488_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1485: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1488_wire_constant & nCOUNTER_1498_1489_buffered;
      req <= phi_stmt_1485_req_0 & phi_stmt_1485_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1485",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1485_ack_0,
          idata => idata,
          odata => COUNTER_1485,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1485
    nCOUNTER_1498_1489_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_1498_1489_buf_req_0;
      nCOUNTER_1498_1489_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_1498_1489_buf_req_1;
      nCOUNTER_1498_1489_buf_ack_1<= rack(0);
      nCOUNTER_1498_1489_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_1498_1489_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_1498,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_1498_1489_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1490
    process(RPIPE_timer_req_1492_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_1492_wire(0 downto 0);
      req_1490 <= tmp_var; -- 
    end process;
    do_while_stmt_1483_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1504_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1483_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1483_branch_req_0,
          ack0 => do_while_stmt_1483_branch_ack_0,
          ack1 => do_while_stmt_1483_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1497_inst
    process(COUNTER_1485) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_1485, konst_1496_wire_constant, tmp_var);
      nCOUNTER_1498 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_1492_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_1492_inst_req_0;
      RPIPE_timer_req_1492_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_1492_inst_req_1;
      RPIPE_timer_req_1492_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_1492_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_1500_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_1500_inst_req_0;
      WPIPE_timer_resp_1500_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_1500_inst_req_1;
      WPIPE_timer_resp_1500_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_1490(0);
      data_in <= COUNTER_1485;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(9 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module ct_core
  component ct_core is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(9 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module ct_core
  signal ct_core_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal ct_core_tag_out   : std_logic_vector(1 downto 0);
  signal ct_core_start_req : std_logic;
  signal ct_core_start_ack : std_logic;
  signal ct_core_fin_req   : std_logic;
  signal ct_core_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module ct_core
  ct_core_instance:ct_core-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => ct_core_start_req,
      start_ack => ct_core_start_ack,
      fin_req => ct_core_fin_req,
      fin_ack => ct_core_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(17 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(18 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(17 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(9 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(0 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(18 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => ct_core_tag_in,
      tag_out => ct_core_tag_out-- 
    ); -- 
  -- module will be run forever 
  ct_core_tag_in <= (others => '0');
  ct_core_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ct_core_start_req, start_ack => ct_core_start_ack,  fin_req => ct_core_fin_req,  fin_ack => ct_core_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_1: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_stores => 1,
      addr_width => 10,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
