-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendOutput_CP_26_start: Boolean;
  signal sendOutput_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_43_branch_ack_1 : boolean;
  signal if_stmt_43_branch_ack_0 : boolean;
  signal if_stmt_43_branch_req_0 : boolean;
  signal type_cast_52_inst_req_0 : boolean;
  signal type_cast_52_inst_ack_0 : boolean;
  signal type_cast_52_inst_req_1 : boolean;
  signal type_cast_52_inst_ack_1 : boolean;
  signal array_obj_ref_68_index_offset_req_0 : boolean;
  signal array_obj_ref_68_index_offset_ack_0 : boolean;
  signal array_obj_ref_68_index_offset_req_1 : boolean;
  signal array_obj_ref_68_index_offset_ack_1 : boolean;
  signal addr_of_69_final_reg_req_0 : boolean;
  signal addr_of_69_final_reg_ack_0 : boolean;
  signal addr_of_69_final_reg_req_1 : boolean;
  signal addr_of_69_final_reg_ack_1 : boolean;
  signal ptr_deref_73_load_0_req_0 : boolean;
  signal ptr_deref_73_load_0_ack_0 : boolean;
  signal ptr_deref_73_load_0_req_1 : boolean;
  signal ptr_deref_73_load_0_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_164_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_164_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_164_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_164_inst_ack_1 : boolean;
  signal type_cast_77_inst_req_0 : boolean;
  signal type_cast_77_inst_ack_0 : boolean;
  signal type_cast_77_inst_req_1 : boolean;
  signal type_cast_77_inst_ack_1 : boolean;
  signal type_cast_87_inst_req_0 : boolean;
  signal type_cast_87_inst_ack_0 : boolean;
  signal type_cast_87_inst_req_1 : boolean;
  signal type_cast_87_inst_ack_1 : boolean;
  signal type_cast_97_inst_req_0 : boolean;
  signal type_cast_97_inst_ack_0 : boolean;
  signal type_cast_97_inst_req_1 : boolean;
  signal type_cast_97_inst_ack_1 : boolean;
  signal type_cast_107_inst_req_0 : boolean;
  signal type_cast_107_inst_ack_0 : boolean;
  signal type_cast_107_inst_req_1 : boolean;
  signal type_cast_107_inst_ack_1 : boolean;
  signal type_cast_117_inst_req_0 : boolean;
  signal type_cast_117_inst_ack_0 : boolean;
  signal type_cast_117_inst_req_1 : boolean;
  signal type_cast_117_inst_ack_1 : boolean;
  signal type_cast_127_inst_req_0 : boolean;
  signal type_cast_127_inst_ack_0 : boolean;
  signal type_cast_127_inst_req_1 : boolean;
  signal type_cast_127_inst_ack_1 : boolean;
  signal type_cast_137_inst_req_0 : boolean;
  signal type_cast_137_inst_ack_0 : boolean;
  signal type_cast_137_inst_req_1 : boolean;
  signal type_cast_137_inst_ack_1 : boolean;
  signal type_cast_147_inst_req_0 : boolean;
  signal type_cast_147_inst_ack_0 : boolean;
  signal type_cast_147_inst_req_1 : boolean;
  signal type_cast_147_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_149_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_149_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_149_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_149_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_152_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_152_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_152_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_152_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_155_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_155_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_155_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_155_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_158_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_158_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_158_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_158_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_161_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_161_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_161_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_161_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_167_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_167_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_167_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_167_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_170_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_170_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_170_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_170_inst_ack_1 : boolean;
  signal if_stmt_184_branch_req_0 : boolean;
  signal if_stmt_184_branch_ack_1 : boolean;
  signal if_stmt_184_branch_ack_0 : boolean;
  signal phi_stmt_56_req_1 : boolean;
  signal type_cast_59_inst_req_0 : boolean;
  signal type_cast_59_inst_ack_0 : boolean;
  signal type_cast_59_inst_req_1 : boolean;
  signal type_cast_59_inst_ack_1 : boolean;
  signal phi_stmt_56_req_0 : boolean;
  signal phi_stmt_56_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_26: Block -- control-path 
    signal sendOutput_CP_26_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendOutput_CP_26_elements(0) <= sendOutput_CP_26_start;
    sendOutput_CP_26_symbol <= sendOutput_CP_26_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_23/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/branch_block_stmt_23__entry__
      -- CP-element group 0: 	 branch_block_stmt_23/if_stmt_43_else_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_33_to_assign_stmt_42__entry__
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_33_to_assign_stmt_42__exit__
      -- CP-element group 0: 	 branch_block_stmt_23/if_stmt_43__entry__
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_33_to_assign_stmt_42/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/assign_stmt_33_to_assign_stmt_42/$exit
      -- CP-element group 0: 	 branch_block_stmt_23/if_stmt_43_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/if_stmt_43_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_23/if_stmt_43_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_23/if_stmt_43_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_23/R_cmp68_44_place
      -- CP-element group 0: 	 branch_block_stmt_23/if_stmt_43_if_link/$entry
      -- 
    branch_req_64_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_64_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => if_stmt_43_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	4 
    -- CP-element group 1: 	3 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_43_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_23/merge_stmt_49__exit__
      -- CP-element group 1: 	 branch_block_stmt_23/assign_stmt_53__entry__
      -- CP-element group 1: 	 branch_block_stmt_23/if_stmt_43_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_23/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_23/assign_stmt_53/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_update_start_
      -- CP-element group 1: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_23/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_23/merge_stmt_49_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_23/merge_stmt_49_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_23/merge_stmt_49_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_23/merge_stmt_49_PhiAck/dummy
      -- 
    if_choice_transition_69_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_43_branch_ack_1, ack => sendOutput_CP_26_elements(1)); -- 
    rr_86_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_86_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(1), ack => type_cast_52_inst_req_0); -- 
    cr_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(1), ack => type_cast_52_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_23/if_stmt_43_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_23/if_stmt_43_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_23/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_23/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_23/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_73_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_43_branch_ack_0, ack => sendOutput_CP_26_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_Sample/ra
      -- 
    ra_87_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_0, ack => sendOutput_CP_26_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_53__exit__
      -- CP-element group 4: 	 branch_block_stmt_23/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_53/$exit
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_23/assign_stmt_53/type_cast_52_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_23/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_23/bbx_xnph_forx_xbody_PhiReq/phi_stmt_56/$entry
      -- CP-element group 4: 	 branch_block_stmt_23/bbx_xnph_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/$entry
      -- 
    ca_92_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_1, ack => sendOutput_CP_26_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_final_index_sum_regn_Sample/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_68_index_offset_ack_0, ack => sendOutput_CP_26_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_request/req
      -- 
    ack_126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_68_index_offset_ack_1, ack => sendOutput_CP_26_elements(6)); -- 
    req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(6), ack => addr_of_69_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_request/$exit
      -- CP-element group 7: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_request/ack
      -- 
    ack_136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_69_final_reg_ack_0, ack => sendOutput_CP_26_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Sample/word_access_start/word_0/rr
      -- 
    ack_141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_69_final_reg_ack_1, ack => sendOutput_CP_26_elements(8)); -- 
    rr_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(8), ack => ptr_deref_73_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Sample/word_access_start/word_0/ra
      -- 
    ra_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_73_load_0_ack_0, ack => sendOutput_CP_26_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	21 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	25 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/ptr_deref_73_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/ptr_deref_73_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/ptr_deref_73_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/ptr_deref_73_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_Sample/rr
      -- 
    ca_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_73_load_0_ack_1, ack => sendOutput_CP_26_elements(10)); -- 
    rr_227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_97_inst_req_0); -- 
    rr_241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_107_inst_req_0); -- 
    rr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_117_inst_req_0); -- 
    rr_269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_127_inst_req_0); -- 
    rr_283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_137_inst_req_0); -- 
    rr_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_147_inst_req_0); -- 
    rr_213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_87_inst_req_0); -- 
    rr_199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_77_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_Sample/ra
      -- 
    ra_200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_0, ack => sendOutput_CP_26_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	47 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_Update/ca
      -- 
    ca_205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_77_inst_ack_1, ack => sendOutput_CP_26_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_Sample/ra
      -- 
    ra_214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_87_inst_ack_0, ack => sendOutput_CP_26_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	58 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	44 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_Update/ca
      -- 
    ca_219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_87_inst_ack_1, ack => sendOutput_CP_26_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_Sample/ra
      -- 
    ra_228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_97_inst_ack_0, ack => sendOutput_CP_26_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_Update/ca
      -- 
    ca_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_97_inst_ack_1, ack => sendOutput_CP_26_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_Sample/ra
      -- 
    ra_242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_0, ack => sendOutput_CP_26_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	58 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	38 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_Update/ca
      -- 
    ca_247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_1, ack => sendOutput_CP_26_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_Sample/ra
      -- 
    ra_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_117_inst_ack_0, ack => sendOutput_CP_26_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	58 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	35 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_Update/ca
      -- 
    ca_261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_117_inst_ack_1, ack => sendOutput_CP_26_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	10 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_Sample/ra
      -- 
    ra_270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_0, ack => sendOutput_CP_26_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	58 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	32 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_Update/ca
      -- 
    ca_275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_1, ack => sendOutput_CP_26_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_Sample/ra
      -- 
    ra_284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_137_inst_ack_0, ack => sendOutput_CP_26_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	58 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_Update/ca
      -- 
    ca_289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_137_inst_ack_1, ack => sendOutput_CP_26_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_Sample/ra
      -- 
    ra_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_147_inst_ack_0, ack => sendOutput_CP_26_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_Sample/req
      -- 
    ca_303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_147_inst_ack_1, ack => sendOutput_CP_26_elements(26)); -- 
    req_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(26), ack => WPIPE_zeropad_output_pipe_149_inst_req_0); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_update_start_
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_Update/req
      -- 
    ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_149_inst_ack_0, ack => sendOutput_CP_26_elements(27)); -- 
    req_316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(27), ack => WPIPE_zeropad_output_pipe_149_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_149_Update/ack
      -- 
    ack_317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_149_inst_ack_1, ack => sendOutput_CP_26_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_Sample/req
      -- 
    req_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(29), ack => WPIPE_zeropad_output_pipe_152_inst_req_0); -- 
    sendOutput_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(24) & sendOutput_CP_26_elements(28);
      gj_sendOutput_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_update_start_
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_Update/req
      -- 
    ack_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_152_inst_ack_0, ack => sendOutput_CP_26_elements(30)); -- 
    req_330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(30), ack => WPIPE_zeropad_output_pipe_152_inst_req_1); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_152_Update/ack
      -- 
    ack_331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_152_inst_ack_1, ack => sendOutput_CP_26_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	22 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_Sample/req
      -- 
    req_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(32), ack => WPIPE_zeropad_output_pipe_155_inst_req_0); -- 
    sendOutput_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(22) & sendOutput_CP_26_elements(31);
      gj_sendOutput_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_update_start_
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_Update/req
      -- 
    ack_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_155_inst_ack_0, ack => sendOutput_CP_26_elements(33)); -- 
    req_344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(33), ack => WPIPE_zeropad_output_pipe_155_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_155_Update/ack
      -- 
    ack_345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_155_inst_ack_1, ack => sendOutput_CP_26_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	20 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_Sample/req
      -- 
    req_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(35), ack => WPIPE_zeropad_output_pipe_158_inst_req_0); -- 
    sendOutput_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(20) & sendOutput_CP_26_elements(34);
      gj_sendOutput_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_update_start_
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_Update/req
      -- 
    ack_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_158_inst_ack_0, ack => sendOutput_CP_26_elements(36)); -- 
    req_358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(36), ack => WPIPE_zeropad_output_pipe_158_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_158_Update/ack
      -- 
    ack_359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_158_inst_ack_1, ack => sendOutput_CP_26_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	18 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_Sample/req
      -- 
    req_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(38), ack => WPIPE_zeropad_output_pipe_161_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(18) & sendOutput_CP_26_elements(37);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_update_start_
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_Update/req
      -- 
    ack_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_161_inst_ack_0, ack => sendOutput_CP_26_elements(39)); -- 
    req_372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(39), ack => WPIPE_zeropad_output_pipe_161_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_161_Update/ack
      -- 
    ack_373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_161_inst_ack_1, ack => sendOutput_CP_26_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_Sample/req
      -- CP-element group 41: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_sample_start_
      -- 
    req_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(41), ack => WPIPE_zeropad_output_pipe_164_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(16) & sendOutput_CP_26_elements(40);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_Update/req
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_update_start_
      -- 
    ack_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_164_inst_ack_0, ack => sendOutput_CP_26_elements(42)); -- 
    req_386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(42), ack => WPIPE_zeropad_output_pipe_164_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_164_Update/ack
      -- 
    ack_387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_164_inst_ack_1, ack => sendOutput_CP_26_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	14 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_Sample/req
      -- 
    req_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(44), ack => WPIPE_zeropad_output_pipe_167_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(14) & sendOutput_CP_26_elements(43);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_update_start_
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_Update/req
      -- 
    ack_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_167_inst_ack_0, ack => sendOutput_CP_26_elements(45)); -- 
    req_400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(45), ack => WPIPE_zeropad_output_pipe_167_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_167_Update/ack
      -- 
    ack_401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_167_inst_ack_1, ack => sendOutput_CP_26_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	12 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_Sample/req
      -- 
    req_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(47), ack => WPIPE_zeropad_output_pipe_170_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(12) & sendOutput_CP_26_elements(46);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_update_start_
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_Update/req
      -- 
    ack_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_170_inst_ack_0, ack => sendOutput_CP_26_elements(48)); -- 
    req_414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(48), ack => WPIPE_zeropad_output_pipe_170_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/WPIPE_zeropad_output_pipe_170_Update/ack
      -- 
    ack_415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_170_inst_ack_1, ack => sendOutput_CP_26_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183__exit__
      -- CP-element group 50: 	 branch_block_stmt_23/if_stmt_184__entry__
      -- CP-element group 50: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/$exit
      -- CP-element group 50: 	 branch_block_stmt_23/if_stmt_184_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_23/if_stmt_184_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_23/if_stmt_184_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_23/if_stmt_184_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_23/R_exitcond2_185_place
      -- CP-element group 50: 	 branch_block_stmt_23/if_stmt_184_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_23/if_stmt_184_else_link/$entry
      -- 
    branch_req_423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(50), ack => if_stmt_184_branch_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(5) & sendOutput_CP_26_elements(49);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_23/merge_stmt_190__exit__
      -- CP-element group 51: 	 branch_block_stmt_23/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_23/if_stmt_184_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_23/if_stmt_184_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_23/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_23/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_23/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_23/merge_stmt_190_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_23/merge_stmt_190_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_23/merge_stmt_190_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_23/merge_stmt_190_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_23/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_23/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_184_branch_ack_1, ack => sendOutput_CP_26_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_23/if_stmt_184_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_23/if_stmt_184_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_23/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/$entry
      -- CP-element group 52: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/$entry
      -- CP-element group 52: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/SplitProtocol/Update/cr
      -- 
    else_choice_transition_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_184_branch_ack_0, ack => sendOutput_CP_26_elements(52)); -- 
    rr_476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(52), ack => type_cast_59_inst_req_0); -- 
    cr_481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(52), ack => type_cast_59_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_23/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_23/bbx_xnph_forx_xbody_PhiReq/phi_stmt_56/$exit
      -- CP-element group 53: 	 branch_block_stmt_23/bbx_xnph_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_23/bbx_xnph_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_62_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_23/bbx_xnph_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_req
      -- 
    phi_stmt_56_req_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_56_req_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(53), ack => phi_stmt_56_req_1); -- 
    -- Element group sendOutput_CP_26_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendOutput_CP_26_elements(4), ack => sendOutput_CP_26_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/SplitProtocol/Sample/ra
      -- 
    ra_477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_59_inst_ack_0, ack => sendOutput_CP_26_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/SplitProtocol/Update/ca
      -- 
    ca_482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_59_inst_ack_1, ack => sendOutput_CP_26_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/$exit
      -- CP-element group 56: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/$exit
      -- CP-element group 56: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_sources/type_cast_59/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_23/forx_xbody_forx_xbody_PhiReq/phi_stmt_56/phi_stmt_56_req
      -- 
    phi_stmt_56_req_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_56_req_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(56), ack => phi_stmt_56_req_0); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(54) & sendOutput_CP_26_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	53 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_23/merge_stmt_55_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_23/merge_stmt_55_PhiAck/$entry
      -- 
    sendOutput_CP_26_elements(57) <= OrReduce(sendOutput_CP_26_elements(53) & sendOutput_CP_26_elements(56));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	18 
    -- CP-element group 58: 	20 
    -- CP-element group 58: 	22 
    -- CP-element group 58: 	24 
    -- CP-element group 58: 	26 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	12 
    -- CP-element group 58: 	10 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_23/merge_stmt_55__exit__
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183__entry__
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/array_obj_ref_68_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/addr_of_69_complete/req
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/ptr_deref_73_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_77_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_87_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_97_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_107_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_117_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_127_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_137_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_update_start_
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_23/assign_stmt_70_to_assign_stmt_183/type_cast_147_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_23/merge_stmt_55_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_23/merge_stmt_55_PhiAck/phi_stmt_56_ack
      -- 
    phi_stmt_56_ack_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_56_ack_0, ack => sendOutput_CP_26_elements(58)); -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => array_obj_ref_68_index_offset_req_0); -- 
    req_125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => array_obj_ref_68_index_offset_req_1); -- 
    req_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => addr_of_69_final_reg_req_1); -- 
    cr_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => ptr_deref_73_load_0_req_1); -- 
    cr_204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_77_inst_req_1); -- 
    cr_218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_87_inst_req_1); -- 
    cr_232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_97_inst_req_1); -- 
    cr_246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_107_inst_req_1); -- 
    cr_260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_117_inst_req_1); -- 
    cr_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_127_inst_req_1); -- 
    cr_288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_137_inst_req_1); -- 
    cr_302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_147_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	2 
    -- CP-element group 59: 	51 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_23/$exit
      -- CP-element group 59: 	 branch_block_stmt_23/branch_block_stmt_23__exit__
      -- CP-element group 59: 	 branch_block_stmt_23/merge_stmt_192__exit__
      -- CP-element group 59: 	 branch_block_stmt_23/return__
      -- CP-element group 59: 	 branch_block_stmt_23/merge_stmt_194__exit__
      -- CP-element group 59: 	 branch_block_stmt_23/merge_stmt_192_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_23/merge_stmt_192_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_23/merge_stmt_192_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_23/merge_stmt_192_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_23/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_23/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_23/merge_stmt_194_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_23/merge_stmt_194_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_23/merge_stmt_194_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_23/merge_stmt_194_PhiAck/dummy
      -- 
    sendOutput_CP_26_elements(59) <= OrReduce(sendOutput_CP_26_elements(2) & sendOutput_CP_26_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_31_wire : std_logic_vector(31 downto 0);
    signal R_indvar_67_resized : std_logic_vector(13 downto 0);
    signal R_indvar_67_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_68_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_68_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_68_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_68_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_68_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_68_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_70 : std_logic_vector(31 downto 0);
    signal cmp68_42 : std_logic_vector(0 downto 0);
    signal conv12_88 : std_logic_vector(7 downto 0);
    signal conv18_98 : std_logic_vector(7 downto 0);
    signal conv24_108 : std_logic_vector(7 downto 0);
    signal conv30_118 : std_logic_vector(7 downto 0);
    signal conv36_128 : std_logic_vector(7 downto 0);
    signal conv42_138 : std_logic_vector(7 downto 0);
    signal conv48_148 : std_logic_vector(7 downto 0);
    signal conv_78 : std_logic_vector(7 downto 0);
    signal exitcond2_183 : std_logic_vector(0 downto 0);
    signal indvar_56 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_178 : std_logic_vector(63 downto 0);
    signal ptr_deref_73_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_73_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_73_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_73_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_73_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_94 : std_logic_vector(63 downto 0);
    signal shr21_104 : std_logic_vector(63 downto 0);
    signal shr27_114 : std_logic_vector(63 downto 0);
    signal shr33_124 : std_logic_vector(63 downto 0);
    signal shr39_134 : std_logic_vector(63 downto 0);
    signal shr45_144 : std_logic_vector(63 downto 0);
    signal shr67_33 : std_logic_vector(31 downto 0);
    signal shr9_84 : std_logic_vector(63 downto 0);
    signal tmp1_53 : std_logic_vector(63 downto 0);
    signal tmp4_74 : std_logic_vector(63 downto 0);
    signal type_cast_102_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_112_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_122_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_132_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_142_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_176_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_27_wire : std_logic_vector(31 downto 0);
    signal type_cast_30_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_36_wire : std_logic_vector(31 downto 0);
    signal type_cast_39_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_59_wire : std_logic_vector(63 downto 0);
    signal type_cast_62_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_82_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_92_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_68_constant_part_of_offset <= "00000000000000";
    array_obj_ref_68_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_68_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_68_resized_base_address <= "00000000000000";
    ptr_deref_73_word_offset_0 <= "00000000000000";
    type_cast_102_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_112_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_122_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_132_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_142_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_176_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_30_wire_constant <= "00000000000000000000000000000010";
    type_cast_39_wire_constant <= "00000000000000000000000000000000";
    type_cast_62_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_82_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_92_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    phi_stmt_56: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_59_wire & type_cast_62_wire_constant;
      req <= phi_stmt_56_req_0 & phi_stmt_56_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_56",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_56_ack_0,
          idata => idata,
          odata => indvar_56,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_56
    addr_of_69_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_69_final_reg_req_0;
      addr_of_69_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_69_final_reg_req_1;
      addr_of_69_final_reg_ack_1<= rack(0);
      addr_of_69_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_69_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_68_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_70,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_107_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_107_inst_req_0;
      type_cast_107_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_107_inst_req_1;
      type_cast_107_inst_ack_1<= rack(0);
      type_cast_107_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_107_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_104,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_108,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_117_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_117_inst_req_0;
      type_cast_117_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_117_inst_req_1;
      type_cast_117_inst_ack_1<= rack(0);
      type_cast_117_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_117_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_114,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_118,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_127_inst_req_0;
      type_cast_127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_127_inst_req_1;
      type_cast_127_inst_ack_1<= rack(0);
      type_cast_127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_137_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_137_inst_req_0;
      type_cast_137_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_137_inst_req_1;
      type_cast_137_inst_ack_1<= rack(0);
      type_cast_137_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_137_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_134,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_138,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_147_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_147_inst_req_0;
      type_cast_147_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_147_inst_req_1;
      type_cast_147_inst_ack_1<= rack(0);
      type_cast_147_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_147_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_144,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_148,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_27_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := size_buffer(31 downto 0);
      type_cast_27_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_32_inst
    process(ASHR_i32_i32_31_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_31_wire(31 downto 0);
      shr67_33 <= tmp_var; -- 
    end process;
    -- interlock type_cast_36_inst
    process(shr67_33) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := shr67_33(31 downto 0);
      type_cast_36_wire <= tmp_var; -- 
    end process;
    type_cast_52_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_52_inst_req_0;
      type_cast_52_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_52_inst_req_1;
      type_cast_52_inst_ack_1<= rack(0);
      type_cast_52_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_52_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr67_33,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_53,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_59_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_59_inst_req_0;
      type_cast_59_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_59_inst_req_1;
      type_cast_59_inst_ack_1<= rack(0);
      type_cast_59_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_59_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_178,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_59_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_77_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_77_inst_req_0;
      type_cast_77_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_77_inst_req_1;
      type_cast_77_inst_ack_1<= rack(0);
      type_cast_77_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_77_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_74,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_78,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_87_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_87_inst_req_0;
      type_cast_87_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_87_inst_req_1;
      type_cast_87_inst_ack_1<= rack(0);
      type_cast_87_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_87_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_84,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_88,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_97_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_97_inst_req_0;
      type_cast_97_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_97_inst_req_1;
      type_cast_97_inst_ack_1<= rack(0);
      type_cast_97_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_97_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_94,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_98,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_68_index_1_rename
    process(R_indvar_67_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_67_resized;
      ov(13 downto 0) := iv;
      R_indvar_67_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_68_index_1_resize
    process(indvar_56) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_56;
      ov := iv(13 downto 0);
      R_indvar_67_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_68_root_address_inst
    process(array_obj_ref_68_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_68_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_68_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_73_addr_0
    process(ptr_deref_73_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_73_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_73_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_73_base_resize
    process(arrayidx_70) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_70;
      ov := iv(13 downto 0);
      ptr_deref_73_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_73_gather_scatter
    process(ptr_deref_73_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_73_data_0;
      ov(63 downto 0) := iv;
      tmp4_74 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_73_root_address_inst
    process(ptr_deref_73_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_73_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_73_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_184_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_183;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_184_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_184_branch_req_0,
          ack0 => if_stmt_184_branch_ack_0,
          ack1 => if_stmt_184_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_43_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp68_42;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_43_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_43_branch_req_0,
          ack0 => if_stmt_43_branch_ack_0,
          ack1 => if_stmt_43_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_177_inst
    process(indvar_56) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_56, type_cast_176_wire_constant, tmp_var);
      indvarx_xnext_178 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_31_inst
    process(type_cast_27_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_27_wire, type_cast_30_wire_constant, tmp_var);
      ASHR_i32_i32_31_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_182_inst
    process(indvarx_xnext_178, tmp1_53) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_178, tmp1_53, tmp_var);
      exitcond2_183 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_103_inst
    process(tmp4_74) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_74, type_cast_102_wire_constant, tmp_var);
      shr21_104 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_113_inst
    process(tmp4_74) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_74, type_cast_112_wire_constant, tmp_var);
      shr27_114 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_123_inst
    process(tmp4_74) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_74, type_cast_122_wire_constant, tmp_var);
      shr33_124 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_133_inst
    process(tmp4_74) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_74, type_cast_132_wire_constant, tmp_var);
      shr39_134 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_143_inst
    process(tmp4_74) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_74, type_cast_142_wire_constant, tmp_var);
      shr45_144 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_83_inst
    process(tmp4_74) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_74, type_cast_82_wire_constant, tmp_var);
      shr9_84 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_93_inst
    process(tmp4_74) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_74, type_cast_92_wire_constant, tmp_var);
      shr15_94 <= tmp_var; --
    end process;
    -- binary operator SGT_i32_u1_40_inst
    process(type_cast_36_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(type_cast_36_wire, type_cast_39_wire_constant, tmp_var);
      cmp68_42 <= tmp_var; --
    end process;
    -- shared split operator group (11) : array_obj_ref_68_index_offset 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_67_scaled;
      array_obj_ref_68_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_68_index_offset_req_0;
      array_obj_ref_68_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_68_index_offset_req_1;
      array_obj_ref_68_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_11_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared load operator group (0) : ptr_deref_73_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_73_load_0_req_0;
      ptr_deref_73_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_73_load_0_req_1;
      ptr_deref_73_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_73_word_address_0;
      ptr_deref_73_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 5,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_149_inst WPIPE_zeropad_output_pipe_152_inst WPIPE_zeropad_output_pipe_155_inst WPIPE_zeropad_output_pipe_158_inst WPIPE_zeropad_output_pipe_161_inst WPIPE_zeropad_output_pipe_164_inst WPIPE_zeropad_output_pipe_167_inst WPIPE_zeropad_output_pipe_170_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_149_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_152_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_155_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_158_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_161_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_164_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_167_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_170_inst_req_0;
      WPIPE_zeropad_output_pipe_149_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_152_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_155_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_158_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_161_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_164_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_167_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_170_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_149_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_152_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_155_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_158_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_161_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_164_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_167_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_170_inst_req_1;
      WPIPE_zeropad_output_pipe_149_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_152_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_155_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_158_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_161_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_164_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_167_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_170_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv48_148 & conv42_138 & conv36_128 & conv30_118 & conv24_108 & conv18_98 & conv12_88 & conv_78;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(3 downto 0);
    zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_data : out  std_logic_vector(31 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D;
architecture zeropad3D_arch of zeropad3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_CP_676_start: Boolean;
  signal zeropad3D_CP_676_symbol: Boolean;
  -- volatile/operator module components. 
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_685_inst_ack_0 : boolean;
  signal type_cast_762_inst_ack_0 : boolean;
  signal type_cast_722_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_475_inst_ack_1 : boolean;
  signal addr_of_1286_final_reg_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_439_inst_req_0 : boolean;
  signal type_cast_520_inst_ack_1 : boolean;
  signal type_cast_685_inst_req_1 : boolean;
  signal type_cast_528_inst_ack_0 : boolean;
  signal type_cast_461_inst_req_1 : boolean;
  signal type_cast_1345_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_439_inst_ack_0 : boolean;
  signal addr_of_1286_final_reg_req_0 : boolean;
  signal type_cast_461_inst_ack_1 : boolean;
  signal type_cast_685_inst_req_0 : boolean;
  signal type_cast_762_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_475_inst_ack_0 : boolean;
  signal LOAD_pad_512_load_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_457_inst_ack_0 : boolean;
  signal LOAD_pad_512_load_0_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_457_inst_req_0 : boolean;
  signal ptr_deref_487_store_0_ack_1 : boolean;
  signal if_stmt_501_branch_req_0 : boolean;
  signal if_stmt_675_branch_req_0 : boolean;
  signal type_cast_524_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_475_inst_req_0 : boolean;
  signal ptr_deref_1289_store_0_req_0 : boolean;
  signal type_cast_1412_inst_req_0 : boolean;
  signal addr_of_769_final_reg_req_0 : boolean;
  signal type_cast_528_inst_req_1 : boolean;
  signal type_cast_722_inst_req_0 : boolean;
  signal type_cast_762_inst_req_1 : boolean;
  signal type_cast_461_inst_ack_0 : boolean;
  signal type_cast_528_inst_ack_1 : boolean;
  signal if_stmt_501_branch_ack_0 : boolean;
  signal type_cast_685_inst_ack_1 : boolean;
  signal type_cast_461_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_475_inst_req_1 : boolean;
  signal type_cast_520_inst_req_1 : boolean;
  signal addr_of_1286_final_reg_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_439_inst_req_1 : boolean;
  signal addr_of_1261_final_reg_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_439_inst_ack_1 : boolean;
  signal ptr_deref_2077_load_0_req_0 : boolean;
  signal type_cast_528_inst_req_0 : boolean;
  signal if_stmt_501_branch_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_457_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_457_inst_ack_1 : boolean;
  signal ptr_deref_487_store_0_req_1 : boolean;
  signal type_cast_425_inst_ack_1 : boolean;
  signal type_cast_443_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_225_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_225_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_225_inst_req_1 : boolean;
  signal type_cast_1345_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_225_inst_ack_1 : boolean;
  signal type_cast_520_inst_ack_0 : boolean;
  signal type_cast_425_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_228_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_228_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_228_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_228_inst_ack_1 : boolean;
  signal if_stmt_712_branch_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_231_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_231_inst_ack_0 : boolean;
  signal type_cast_727_inst_ack_1 : boolean;
  signal type_cast_1509_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_231_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_231_inst_ack_1 : boolean;
  signal addr_of_769_final_reg_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_234_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_234_inst_ack_0 : boolean;
  signal addr_of_769_final_reg_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_234_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_234_inst_ack_1 : boolean;
  signal if_stmt_712_branch_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_237_inst_req_0 : boolean;
  signal type_cast_648_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_237_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_237_inst_req_1 : boolean;
  signal type_cast_648_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_237_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_240_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_240_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_240_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_240_inst_ack_1 : boolean;
  signal type_cast_520_inst_req_0 : boolean;
  signal type_cast_727_inst_req_1 : boolean;
  signal addr_of_1286_final_reg_ack_1 : boolean;
  signal type_cast_648_inst_ack_0 : boolean;
  signal type_cast_648_inst_req_0 : boolean;
  signal ptr_deref_487_store_0_ack_0 : boolean;
  signal addr_of_769_final_reg_ack_0 : boolean;
  signal STORE_pad_242_store_0_req_0 : boolean;
  signal STORE_pad_242_store_0_ack_0 : boolean;
  signal type_cast_443_inst_req_1 : boolean;
  signal ptr_deref_487_store_0_req_0 : boolean;
  signal STORE_pad_242_store_0_req_1 : boolean;
  signal STORE_pad_242_store_0_ack_1 : boolean;
  signal ptr_deref_772_store_0_req_1 : boolean;
  signal array_obj_ref_1285_index_offset_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_246_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_246_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_246_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_246_inst_ack_1 : boolean;
  signal if_stmt_712_branch_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_249_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_249_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_249_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_249_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_252_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_252_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_252_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_252_inst_ack_1 : boolean;
  signal type_cast_1509_inst_req_1 : boolean;
  signal type_cast_256_inst_req_0 : boolean;
  signal type_cast_256_inst_ack_0 : boolean;
  signal type_cast_256_inst_req_1 : boolean;
  signal type_cast_256_inst_ack_1 : boolean;
  signal type_cast_727_inst_ack_0 : boolean;
  signal type_cast_260_inst_req_0 : boolean;
  signal type_cast_577_inst_ack_1 : boolean;
  signal type_cast_260_inst_ack_0 : boolean;
  signal type_cast_260_inst_req_1 : boolean;
  signal type_cast_577_inst_req_1 : boolean;
  signal type_cast_260_inst_ack_1 : boolean;
  signal type_cast_727_inst_req_0 : boolean;
  signal type_cast_264_inst_req_0 : boolean;
  signal type_cast_264_inst_ack_0 : boolean;
  signal type_cast_264_inst_req_1 : boolean;
  signal type_cast_264_inst_ack_1 : boolean;
  signal type_cast_516_inst_ack_1 : boolean;
  signal if_stmt_288_branch_req_0 : boolean;
  signal type_cast_516_inst_req_1 : boolean;
  signal type_cast_524_inst_ack_1 : boolean;
  signal type_cast_443_inst_ack_0 : boolean;
  signal if_stmt_288_branch_ack_1 : boolean;
  signal type_cast_524_inst_req_1 : boolean;
  signal type_cast_443_inst_req_0 : boolean;
  signal if_stmt_288_branch_ack_0 : boolean;
  signal type_cast_1345_inst_req_1 : boolean;
  signal type_cast_297_inst_req_0 : boolean;
  signal type_cast_577_inst_ack_0 : boolean;
  signal type_cast_297_inst_ack_0 : boolean;
  signal type_cast_297_inst_req_1 : boolean;
  signal type_cast_577_inst_req_0 : boolean;
  signal type_cast_297_inst_ack_1 : boolean;
  signal if_stmt_1536_branch_req_0 : boolean;
  signal type_cast_301_inst_req_0 : boolean;
  signal type_cast_301_inst_ack_0 : boolean;
  signal type_cast_301_inst_req_1 : boolean;
  signal type_cast_301_inst_ack_1 : boolean;
  signal addr_of_1261_final_reg_ack_0 : boolean;
  signal type_cast_310_inst_req_0 : boolean;
  signal type_cast_310_inst_ack_0 : boolean;
  signal type_cast_310_inst_req_1 : boolean;
  signal type_cast_310_inst_ack_1 : boolean;
  signal type_cast_516_inst_ack_0 : boolean;
  signal if_stmt_675_branch_ack_0 : boolean;
  signal type_cast_516_inst_req_0 : boolean;
  signal type_cast_524_inst_ack_0 : boolean;
  signal LOAD_pad_1408_load_0_req_1 : boolean;
  signal array_obj_ref_350_index_offset_req_0 : boolean;
  signal array_obj_ref_350_index_offset_ack_0 : boolean;
  signal array_obj_ref_350_index_offset_req_1 : boolean;
  signal array_obj_ref_350_index_offset_ack_1 : boolean;
  signal type_cast_541_inst_ack_1 : boolean;
  signal type_cast_479_inst_ack_1 : boolean;
  signal type_cast_541_inst_req_1 : boolean;
  signal addr_of_351_final_reg_req_0 : boolean;
  signal addr_of_351_final_reg_ack_0 : boolean;
  signal addr_of_351_final_reg_req_1 : boolean;
  signal addr_of_351_final_reg_ack_1 : boolean;
  signal array_obj_ref_768_index_offset_ack_1 : boolean;
  signal ptr_deref_772_store_0_ack_0 : boolean;
  signal LOAD_pad_1408_load_0_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_354_inst_req_0 : boolean;
  signal type_cast_541_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_354_inst_ack_0 : boolean;
  signal type_cast_479_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_354_inst_req_1 : boolean;
  signal type_cast_541_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_354_inst_ack_1 : boolean;
  signal ptr_deref_1289_store_0_ack_0 : boolean;
  signal type_cast_358_inst_req_0 : boolean;
  signal type_cast_358_inst_ack_0 : boolean;
  signal type_cast_358_inst_req_1 : boolean;
  signal type_cast_358_inst_ack_1 : boolean;
  signal array_obj_ref_768_index_offset_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_367_inst_ack_1 : boolean;
  signal if_stmt_675_branch_ack_1 : boolean;
  signal type_cast_722_inst_ack_1 : boolean;
  signal type_cast_371_inst_req_0 : boolean;
  signal type_cast_371_inst_ack_0 : boolean;
  signal type_cast_371_inst_req_1 : boolean;
  signal type_cast_371_inst_ack_1 : boolean;
  signal ptr_deref_772_store_0_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_385_inst_req_0 : boolean;
  signal type_cast_537_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_385_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_385_inst_req_1 : boolean;
  signal type_cast_537_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_385_inst_ack_1 : boolean;
  signal type_cast_389_inst_req_0 : boolean;
  signal type_cast_389_inst_ack_0 : boolean;
  signal type_cast_389_inst_req_1 : boolean;
  signal type_cast_389_inst_ack_1 : boolean;
  signal array_obj_ref_768_index_offset_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_403_inst_req_0 : boolean;
  signal type_cast_537_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_403_inst_ack_0 : boolean;
  signal type_cast_479_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_403_inst_req_1 : boolean;
  signal type_cast_537_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_403_inst_ack_1 : boolean;
  signal type_cast_1509_inst_ack_1 : boolean;
  signal LOAD_pad_512_load_0_ack_1 : boolean;
  signal type_cast_722_inst_req_1 : boolean;
  signal type_cast_407_inst_req_0 : boolean;
  signal type_cast_407_inst_ack_0 : boolean;
  signal type_cast_407_inst_req_1 : boolean;
  signal type_cast_407_inst_ack_1 : boolean;
  signal ptr_deref_772_store_0_ack_1 : boolean;
  signal array_obj_ref_768_index_offset_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_421_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_421_inst_ack_0 : boolean;
  signal type_cast_479_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_421_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_421_inst_ack_1 : boolean;
  signal type_cast_762_inst_ack_1 : boolean;
  signal LOAD_pad_512_load_0_req_1 : boolean;
  signal type_cast_425_inst_req_0 : boolean;
  signal type_cast_1345_inst_ack_1 : boolean;
  signal type_cast_425_inst_ack_0 : boolean;
  signal addr_of_1261_final_reg_req_0 : boolean;
  signal type_cast_1336_inst_ack_1 : boolean;
  signal type_cast_1336_inst_req_1 : boolean;
  signal type_cast_781_inst_req_0 : boolean;
  signal type_cast_781_inst_ack_0 : boolean;
  signal if_stmt_1499_branch_ack_0 : boolean;
  signal type_cast_781_inst_req_1 : boolean;
  signal type_cast_781_inst_ack_1 : boolean;
  signal array_obj_ref_2097_index_offset_ack_1 : boolean;
  signal type_cast_1399_inst_ack_1 : boolean;
  signal array_obj_ref_1285_index_offset_req_1 : boolean;
  signal type_cast_845_inst_req_0 : boolean;
  signal type_cast_1336_inst_ack_0 : boolean;
  signal type_cast_845_inst_ack_0 : boolean;
  signal if_stmt_1499_branch_ack_1 : boolean;
  signal type_cast_845_inst_req_1 : boolean;
  signal type_cast_1336_inst_req_0 : boolean;
  signal type_cast_845_inst_ack_1 : boolean;
  signal type_cast_1399_inst_req_1 : boolean;
  signal type_cast_1399_inst_ack_0 : boolean;
  signal type_cast_1399_inst_req_0 : boolean;
  signal array_obj_ref_1285_index_offset_ack_0 : boolean;
  signal array_obj_ref_1285_index_offset_req_0 : boolean;
  signal ptr_deref_2077_load_0_ack_0 : boolean;
  signal array_obj_ref_851_index_offset_req_0 : boolean;
  signal array_obj_ref_851_index_offset_ack_0 : boolean;
  signal array_obj_ref_851_index_offset_req_1 : boolean;
  signal array_obj_ref_851_index_offset_ack_1 : boolean;
  signal type_cast_1509_inst_req_0 : boolean;
  signal if_stmt_1499_branch_req_0 : boolean;
  signal addr_of_852_final_reg_req_0 : boolean;
  signal addr_of_852_final_reg_ack_0 : boolean;
  signal addr_of_852_final_reg_req_1 : boolean;
  signal addr_of_852_final_reg_ack_1 : boolean;
  signal ptr_deref_1265_load_0_ack_0 : boolean;
  signal ptr_deref_1265_load_0_req_0 : boolean;
  signal ptr_deref_856_load_0_req_0 : boolean;
  signal ptr_deref_856_load_0_ack_0 : boolean;
  signal ptr_deref_856_load_0_req_1 : boolean;
  signal ptr_deref_856_load_0_ack_1 : boolean;
  signal if_stmt_1312_branch_ack_0 : boolean;
  signal array_obj_ref_1260_index_offset_ack_1 : boolean;
  signal array_obj_ref_1260_index_offset_req_1 : boolean;
  signal if_stmt_1368_branch_ack_0 : boolean;
  signal type_cast_870_inst_req_0 : boolean;
  signal type_cast_870_inst_ack_0 : boolean;
  signal type_cast_870_inst_req_1 : boolean;
  signal type_cast_870_inst_ack_1 : boolean;
  signal if_stmt_1368_branch_ack_1 : boolean;
  signal if_stmt_1368_branch_req_0 : boolean;
  signal array_obj_ref_876_index_offset_req_0 : boolean;
  signal if_stmt_1312_branch_ack_1 : boolean;
  signal array_obj_ref_876_index_offset_ack_0 : boolean;
  signal array_obj_ref_876_index_offset_req_1 : boolean;
  signal array_obj_ref_876_index_offset_ack_1 : boolean;
  signal if_stmt_1312_branch_req_0 : boolean;
  signal type_cast_1472_inst_ack_1 : boolean;
  signal addr_of_877_final_reg_req_0 : boolean;
  signal addr_of_877_final_reg_ack_0 : boolean;
  signal type_cast_1472_inst_req_1 : boolean;
  signal addr_of_877_final_reg_req_1 : boolean;
  signal addr_of_877_final_reg_ack_1 : boolean;
  signal type_cast_1361_inst_ack_1 : boolean;
  signal type_cast_1361_inst_req_1 : boolean;
  signal type_cast_1297_inst_ack_1 : boolean;
  signal ptr_deref_880_store_0_req_0 : boolean;
  signal ptr_deref_880_store_0_ack_0 : boolean;
  signal ptr_deref_880_store_0_req_1 : boolean;
  signal ptr_deref_880_store_0_ack_1 : boolean;
  signal type_cast_1279_inst_ack_1 : boolean;
  signal type_cast_1361_inst_ack_0 : boolean;
  signal type_cast_888_inst_req_0 : boolean;
  signal type_cast_1297_inst_req_1 : boolean;
  signal type_cast_888_inst_ack_0 : boolean;
  signal type_cast_1472_inst_ack_0 : boolean;
  signal type_cast_888_inst_req_1 : boolean;
  signal type_cast_888_inst_ack_1 : boolean;
  signal LOAD_pad_1408_load_0_ack_0 : boolean;
  signal type_cast_1472_inst_req_0 : boolean;
  signal array_obj_ref_1260_index_offset_ack_0 : boolean;
  signal if_stmt_903_branch_req_0 : boolean;
  signal type_cast_1279_inst_req_1 : boolean;
  signal array_obj_ref_1260_index_offset_req_0 : boolean;
  signal if_stmt_903_branch_ack_1 : boolean;
  signal if_stmt_903_branch_ack_0 : boolean;
  signal type_cast_1297_inst_ack_0 : boolean;
  signal type_cast_927_inst_req_0 : boolean;
  signal type_cast_1297_inst_req_0 : boolean;
  signal type_cast_927_inst_ack_0 : boolean;
  signal type_cast_927_inst_req_1 : boolean;
  signal type_cast_927_inst_ack_1 : boolean;
  signal type_cast_1361_inst_req_0 : boolean;
  signal type_cast_1279_inst_ack_0 : boolean;
  signal LOAD_pad_1408_load_0_req_0 : boolean;
  signal type_cast_936_inst_req_0 : boolean;
  signal type_cast_936_inst_ack_0 : boolean;
  signal type_cast_936_inst_req_1 : boolean;
  signal type_cast_936_inst_ack_1 : boolean;
  signal type_cast_1279_inst_req_0 : boolean;
  signal type_cast_953_inst_req_0 : boolean;
  signal type_cast_953_inst_ack_0 : boolean;
  signal type_cast_953_inst_req_1 : boolean;
  signal type_cast_953_inst_ack_1 : boolean;
  signal type_cast_1412_inst_ack_0 : boolean;
  signal type_cast_1412_inst_ack_1 : boolean;
  signal if_stmt_960_branch_req_0 : boolean;
  signal if_stmt_960_branch_ack_1 : boolean;
  signal if_stmt_960_branch_ack_0 : boolean;
  signal type_cast_1412_inst_req_1 : boolean;
  signal type_cast_991_inst_req_0 : boolean;
  signal ptr_deref_1289_store_0_ack_1 : boolean;
  signal type_cast_991_inst_ack_0 : boolean;
  signal type_cast_991_inst_req_1 : boolean;
  signal ptr_deref_1289_store_0_req_1 : boolean;
  signal type_cast_991_inst_ack_1 : boolean;
  signal addr_of_1261_final_reg_ack_1 : boolean;
  signal LOAD_pad_1000_load_0_req_0 : boolean;
  signal LOAD_pad_1000_load_0_ack_0 : boolean;
  signal LOAD_pad_1000_load_0_req_1 : boolean;
  signal ptr_deref_1265_load_0_ack_1 : boolean;
  signal LOAD_pad_1000_load_0_ack_1 : boolean;
  signal ptr_deref_1265_load_0_req_1 : boolean;
  signal type_cast_2066_inst_req_1 : boolean;
  signal type_cast_2066_inst_ack_1 : boolean;
  signal type_cast_1004_inst_req_0 : boolean;
  signal type_cast_1004_inst_ack_0 : boolean;
  signal type_cast_1004_inst_req_1 : boolean;
  signal type_cast_1004_inst_ack_1 : boolean;
  signal addr_of_2098_final_reg_req_0 : boolean;
  signal type_cast_1058_inst_req_0 : boolean;
  signal addr_of_2098_final_reg_ack_0 : boolean;
  signal type_cast_1058_inst_ack_0 : boolean;
  signal type_cast_1058_inst_req_1 : boolean;
  signal type_cast_1058_inst_ack_1 : boolean;
  signal if_stmt_1085_branch_req_0 : boolean;
  signal if_stmt_1085_branch_ack_1 : boolean;
  signal if_stmt_1085_branch_ack_0 : boolean;
  signal type_cast_1095_inst_req_0 : boolean;
  signal type_cast_1095_inst_ack_0 : boolean;
  signal type_cast_2109_inst_req_0 : boolean;
  signal type_cast_1095_inst_req_1 : boolean;
  signal type_cast_1095_inst_ack_1 : boolean;
  signal if_stmt_2124_branch_ack_0 : boolean;
  signal ptr_deref_1993_store_0_req_1 : boolean;
  signal ptr_deref_1993_store_0_ack_1 : boolean;
  signal if_stmt_1122_branch_req_0 : boolean;
  signal if_stmt_1122_branch_ack_1 : boolean;
  signal if_stmt_1122_branch_ack_0 : boolean;
  signal type_cast_2109_inst_ack_0 : boolean;
  signal type_cast_1132_inst_req_0 : boolean;
  signal type_cast_1132_inst_ack_0 : boolean;
  signal type_cast_1132_inst_req_1 : boolean;
  signal type_cast_1132_inst_ack_1 : boolean;
  signal type_cast_1137_inst_req_0 : boolean;
  signal type_cast_1137_inst_ack_0 : boolean;
  signal type_cast_1137_inst_req_1 : boolean;
  signal type_cast_1137_inst_ack_1 : boolean;
  signal type_cast_1171_inst_req_0 : boolean;
  signal type_cast_1171_inst_ack_0 : boolean;
  signal type_cast_1171_inst_req_1 : boolean;
  signal type_cast_1171_inst_ack_1 : boolean;
  signal ptr_deref_2077_load_0_req_1 : boolean;
  signal if_stmt_2124_branch_ack_1 : boolean;
  signal array_obj_ref_1177_index_offset_req_0 : boolean;
  signal array_obj_ref_1177_index_offset_ack_0 : boolean;
  signal array_obj_ref_1177_index_offset_req_1 : boolean;
  signal array_obj_ref_1177_index_offset_ack_1 : boolean;
  signal addr_of_1178_final_reg_req_0 : boolean;
  signal addr_of_1178_final_reg_ack_0 : boolean;
  signal addr_of_1178_final_reg_req_1 : boolean;
  signal addr_of_1178_final_reg_ack_1 : boolean;
  signal ptr_deref_1181_store_0_req_0 : boolean;
  signal ptr_deref_1181_store_0_ack_0 : boolean;
  signal ptr_deref_1181_store_0_req_1 : boolean;
  signal ptr_deref_1181_store_0_ack_1 : boolean;
  signal type_cast_1190_inst_req_0 : boolean;
  signal type_cast_1190_inst_ack_0 : boolean;
  signal type_cast_1190_inst_req_1 : boolean;
  signal type_cast_1190_inst_ack_1 : boolean;
  signal type_cast_1254_inst_req_0 : boolean;
  signal type_cast_1254_inst_ack_0 : boolean;
  signal type_cast_1254_inst_req_1 : boolean;
  signal type_cast_1254_inst_ack_1 : boolean;
  signal array_obj_ref_2097_index_offset_req_1 : boolean;
  signal if_stmt_1536_branch_ack_1 : boolean;
  signal if_stmt_1536_branch_ack_0 : boolean;
  signal type_cast_1546_inst_req_0 : boolean;
  signal array_obj_ref_2097_index_offset_ack_0 : boolean;
  signal type_cast_1546_inst_ack_0 : boolean;
  signal type_cast_1546_inst_req_1 : boolean;
  signal array_obj_ref_2097_index_offset_req_0 : boolean;
  signal type_cast_1546_inst_ack_1 : boolean;
  signal ptr_deref_2101_store_0_ack_1 : boolean;
  signal type_cast_1551_inst_req_0 : boolean;
  signal type_cast_1551_inst_ack_0 : boolean;
  signal ptr_deref_2101_store_0_req_1 : boolean;
  signal type_cast_1551_inst_req_1 : boolean;
  signal type_cast_1551_inst_ack_1 : boolean;
  signal type_cast_2066_inst_ack_0 : boolean;
  signal type_cast_2066_inst_req_0 : boolean;
  signal type_cast_1585_inst_req_0 : boolean;
  signal type_cast_1585_inst_ack_0 : boolean;
  signal type_cast_1585_inst_req_1 : boolean;
  signal type_cast_1585_inst_ack_1 : boolean;
  signal if_stmt_2124_branch_req_0 : boolean;
  signal array_obj_ref_1591_index_offset_req_0 : boolean;
  signal array_obj_ref_1591_index_offset_ack_0 : boolean;
  signal array_obj_ref_1591_index_offset_req_1 : boolean;
  signal array_obj_ref_1591_index_offset_ack_1 : boolean;
  signal addr_of_1592_final_reg_req_0 : boolean;
  signal addr_of_1592_final_reg_ack_0 : boolean;
  signal addr_of_1592_final_reg_req_1 : boolean;
  signal addr_of_1592_final_reg_ack_1 : boolean;
  signal addr_of_2073_final_reg_ack_1 : boolean;
  signal type_cast_2002_inst_ack_1 : boolean;
  signal addr_of_2073_final_reg_req_1 : boolean;
  signal ptr_deref_1993_store_0_ack_0 : boolean;
  signal ptr_deref_1993_store_0_req_0 : boolean;
  signal ptr_deref_1595_store_0_req_0 : boolean;
  signal ptr_deref_1595_store_0_ack_0 : boolean;
  signal ptr_deref_1595_store_0_req_1 : boolean;
  signal addr_of_2073_final_reg_ack_0 : boolean;
  signal ptr_deref_1595_store_0_ack_1 : boolean;
  signal type_cast_2002_inst_req_1 : boolean;
  signal addr_of_2073_final_reg_req_0 : boolean;
  signal type_cast_1604_inst_req_0 : boolean;
  signal type_cast_1604_inst_ack_0 : boolean;
  signal ptr_deref_2077_load_0_ack_1 : boolean;
  signal ptr_deref_2101_store_0_ack_0 : boolean;
  signal type_cast_1604_inst_req_1 : boolean;
  signal type_cast_1604_inst_ack_1 : boolean;
  signal type_cast_2002_inst_ack_0 : boolean;
  signal ptr_deref_2101_store_0_req_0 : boolean;
  signal type_cast_1668_inst_req_0 : boolean;
  signal type_cast_1668_inst_ack_0 : boolean;
  signal type_cast_1668_inst_req_1 : boolean;
  signal type_cast_2091_inst_ack_1 : boolean;
  signal type_cast_1668_inst_ack_1 : boolean;
  signal type_cast_2002_inst_req_0 : boolean;
  signal array_obj_ref_2072_index_offset_ack_1 : boolean;
  signal array_obj_ref_2072_index_offset_req_1 : boolean;
  signal array_obj_ref_2072_index_offset_ack_0 : boolean;
  signal array_obj_ref_2072_index_offset_req_0 : boolean;
  signal array_obj_ref_1674_index_offset_req_0 : boolean;
  signal type_cast_2091_inst_req_1 : boolean;
  signal array_obj_ref_1674_index_offset_ack_0 : boolean;
  signal array_obj_ref_1674_index_offset_req_1 : boolean;
  signal array_obj_ref_1674_index_offset_ack_1 : boolean;
  signal type_cast_2109_inst_ack_1 : boolean;
  signal type_cast_2109_inst_req_1 : boolean;
  signal type_cast_2091_inst_ack_0 : boolean;
  signal addr_of_1675_final_reg_req_0 : boolean;
  signal type_cast_2091_inst_req_0 : boolean;
  signal addr_of_1675_final_reg_ack_0 : boolean;
  signal addr_of_1675_final_reg_req_1 : boolean;
  signal addr_of_1675_final_reg_ack_1 : boolean;
  signal addr_of_2098_final_reg_ack_1 : boolean;
  signal addr_of_2098_final_reg_req_1 : boolean;
  signal addr_of_2804_final_reg_req_1 : boolean;
  signal ptr_deref_1679_load_0_req_0 : boolean;
  signal ptr_deref_1679_load_0_ack_0 : boolean;
  signal ptr_deref_1679_load_0_req_1 : boolean;
  signal addr_of_2804_final_reg_ack_1 : boolean;
  signal ptr_deref_1679_load_0_ack_1 : boolean;
  signal type_cast_2763_inst_req_1 : boolean;
  signal type_cast_1693_inst_req_0 : boolean;
  signal type_cast_1693_inst_ack_0 : boolean;
  signal type_cast_2763_inst_ack_1 : boolean;
  signal type_cast_1693_inst_req_1 : boolean;
  signal type_cast_1693_inst_ack_1 : boolean;
  signal type_cast_2816_inst_ack_0 : boolean;
  signal type_cast_2816_inst_ack_1 : boolean;
  signal array_obj_ref_1699_index_offset_req_0 : boolean;
  signal array_obj_ref_1699_index_offset_ack_0 : boolean;
  signal array_obj_ref_1699_index_offset_req_1 : boolean;
  signal array_obj_ref_1699_index_offset_ack_1 : boolean;
  signal type_cast_2880_inst_req_0 : boolean;
  signal ptr_deref_2807_store_0_req_1 : boolean;
  signal addr_of_1700_final_reg_req_0 : boolean;
  signal ptr_deref_2807_store_0_ack_1 : boolean;
  signal addr_of_1700_final_reg_ack_0 : boolean;
  signal addr_of_1700_final_reg_req_1 : boolean;
  signal addr_of_1700_final_reg_ack_1 : boolean;
  signal array_obj_ref_2803_index_offset_req_0 : boolean;
  signal ptr_deref_1703_store_0_req_0 : boolean;
  signal ptr_deref_1703_store_0_ack_0 : boolean;
  signal ptr_deref_1703_store_0_req_1 : boolean;
  signal array_obj_ref_2803_index_offset_ack_0 : boolean;
  signal ptr_deref_1703_store_0_ack_1 : boolean;
  signal type_cast_1711_inst_req_0 : boolean;
  signal type_cast_1711_inst_ack_0 : boolean;
  signal type_cast_1711_inst_req_1 : boolean;
  signal type_cast_1711_inst_ack_1 : boolean;
  signal array_obj_ref_2803_index_offset_req_1 : boolean;
  signal array_obj_ref_2803_index_offset_ack_1 : boolean;
  signal if_stmt_1726_branch_req_0 : boolean;
  signal if_stmt_1726_branch_ack_1 : boolean;
  signal if_stmt_1726_branch_ack_0 : boolean;
  signal type_cast_1750_inst_req_0 : boolean;
  signal type_cast_1750_inst_ack_0 : boolean;
  signal type_cast_1750_inst_req_1 : boolean;
  signal type_cast_1750_inst_ack_1 : boolean;
  signal type_cast_1759_inst_req_0 : boolean;
  signal type_cast_1759_inst_ack_0 : boolean;
  signal type_cast_2797_inst_req_0 : boolean;
  signal type_cast_2797_inst_ack_0 : boolean;
  signal type_cast_1759_inst_req_1 : boolean;
  signal type_cast_1759_inst_ack_1 : boolean;
  signal addr_of_2804_final_reg_req_0 : boolean;
  signal type_cast_2816_inst_req_1 : boolean;
  signal type_cast_1776_inst_req_0 : boolean;
  signal type_cast_1776_inst_ack_0 : boolean;
  signal type_cast_1776_inst_req_1 : boolean;
  signal type_cast_1776_inst_ack_1 : boolean;
  signal if_stmt_1783_branch_req_0 : boolean;
  signal if_stmt_1783_branch_ack_1 : boolean;
  signal if_stmt_1783_branch_ack_0 : boolean;
  signal LOAD_pad_1813_load_0_req_0 : boolean;
  signal LOAD_pad_1813_load_0_ack_0 : boolean;
  signal LOAD_pad_1813_load_0_req_1 : boolean;
  signal LOAD_pad_1813_load_0_ack_1 : boolean;
  signal type_cast_1817_inst_req_0 : boolean;
  signal type_cast_1817_inst_ack_0 : boolean;
  signal type_cast_1817_inst_req_1 : boolean;
  signal type_cast_1817_inst_ack_1 : boolean;
  signal type_cast_1870_inst_req_0 : boolean;
  signal type_cast_1870_inst_ack_0 : boolean;
  signal type_cast_1870_inst_req_1 : boolean;
  signal type_cast_1870_inst_ack_1 : boolean;
  signal if_stmt_1897_branch_req_0 : boolean;
  signal if_stmt_1897_branch_ack_1 : boolean;
  signal if_stmt_1897_branch_ack_0 : boolean;
  signal type_cast_1907_inst_req_0 : boolean;
  signal type_cast_1907_inst_ack_0 : boolean;
  signal type_cast_1907_inst_req_1 : boolean;
  signal type_cast_1907_inst_ack_1 : boolean;
  signal if_stmt_1934_branch_req_0 : boolean;
  signal if_stmt_1934_branch_ack_1 : boolean;
  signal if_stmt_1934_branch_ack_0 : boolean;
  signal type_cast_1944_inst_req_0 : boolean;
  signal type_cast_1944_inst_ack_0 : boolean;
  signal type_cast_1944_inst_req_1 : boolean;
  signal type_cast_1944_inst_ack_1 : boolean;
  signal type_cast_1949_inst_req_0 : boolean;
  signal type_cast_1949_inst_ack_0 : boolean;
  signal type_cast_1949_inst_req_1 : boolean;
  signal type_cast_1949_inst_ack_1 : boolean;
  signal type_cast_1983_inst_req_0 : boolean;
  signal type_cast_1983_inst_ack_0 : boolean;
  signal type_cast_1983_inst_req_1 : boolean;
  signal type_cast_1983_inst_ack_1 : boolean;
  signal array_obj_ref_1989_index_offset_req_0 : boolean;
  signal array_obj_ref_1989_index_offset_ack_0 : boolean;
  signal array_obj_ref_1989_index_offset_req_1 : boolean;
  signal array_obj_ref_1989_index_offset_ack_1 : boolean;
  signal addr_of_1990_final_reg_req_0 : boolean;
  signal addr_of_1990_final_reg_ack_0 : boolean;
  signal addr_of_1990_final_reg_req_1 : boolean;
  signal addr_of_1990_final_reg_ack_1 : boolean;
  signal type_cast_2148_inst_req_0 : boolean;
  signal type_cast_2148_inst_ack_0 : boolean;
  signal type_cast_2148_inst_req_1 : boolean;
  signal type_cast_2148_inst_ack_1 : boolean;
  signal type_cast_2157_inst_req_0 : boolean;
  signal type_cast_2157_inst_ack_0 : boolean;
  signal type_cast_2157_inst_req_1 : boolean;
  signal type_cast_2157_inst_ack_1 : boolean;
  signal type_cast_2173_inst_req_0 : boolean;
  signal type_cast_2173_inst_ack_0 : boolean;
  signal type_cast_2173_inst_req_1 : boolean;
  signal type_cast_2173_inst_ack_1 : boolean;
  signal if_stmt_2180_branch_req_0 : boolean;
  signal if_stmt_2180_branch_ack_1 : boolean;
  signal if_stmt_2180_branch_ack_0 : boolean;
  signal LOAD_pad_2216_load_0_req_0 : boolean;
  signal LOAD_pad_2216_load_0_ack_0 : boolean;
  signal LOAD_pad_2216_load_0_req_1 : boolean;
  signal LOAD_pad_2216_load_0_ack_1 : boolean;
  signal type_cast_2220_inst_req_0 : boolean;
  signal type_cast_2220_inst_ack_0 : boolean;
  signal type_cast_2220_inst_req_1 : boolean;
  signal type_cast_2220_inst_ack_1 : boolean;
  signal type_cast_2286_inst_req_0 : boolean;
  signal type_cast_2286_inst_ack_0 : boolean;
  signal type_cast_2286_inst_req_1 : boolean;
  signal ptr_deref_2807_store_0_ack_0 : boolean;
  signal type_cast_2286_inst_ack_1 : boolean;
  signal type_cast_2816_inst_req_0 : boolean;
  signal type_cast_2880_inst_ack_1 : boolean;
  signal if_stmt_2313_branch_req_0 : boolean;
  signal type_cast_2880_inst_req_1 : boolean;
  signal if_stmt_2313_branch_ack_1 : boolean;
  signal type_cast_2763_inst_ack_0 : boolean;
  signal if_stmt_2313_branch_ack_0 : boolean;
  signal ptr_deref_2807_store_0_req_0 : boolean;
  signal type_cast_2323_inst_req_0 : boolean;
  signal type_cast_2323_inst_ack_0 : boolean;
  signal type_cast_2763_inst_req_0 : boolean;
  signal type_cast_2323_inst_req_1 : boolean;
  signal type_cast_2323_inst_ack_1 : boolean;
  signal addr_of_2804_final_reg_ack_0 : boolean;
  signal type_cast_2880_inst_ack_0 : boolean;
  signal type_cast_2797_inst_ack_1 : boolean;
  signal if_stmt_2350_branch_req_0 : boolean;
  signal type_cast_2797_inst_req_1 : boolean;
  signal if_stmt_2350_branch_ack_1 : boolean;
  signal if_stmt_2350_branch_ack_0 : boolean;
  signal type_cast_2360_inst_req_0 : boolean;
  signal type_cast_2360_inst_ack_0 : boolean;
  signal type_cast_2360_inst_req_1 : boolean;
  signal type_cast_2360_inst_ack_1 : boolean;
  signal array_obj_ref_3315_index_offset_ack_1 : boolean;
  signal type_cast_2365_inst_req_0 : boolean;
  signal type_cast_2365_inst_ack_0 : boolean;
  signal type_cast_2365_inst_req_1 : boolean;
  signal type_cast_2365_inst_ack_1 : boolean;
  signal type_cast_2399_inst_req_0 : boolean;
  signal type_cast_2399_inst_ack_0 : boolean;
  signal type_cast_2399_inst_req_1 : boolean;
  signal type_cast_2399_inst_ack_1 : boolean;
  signal type_cast_3366_inst_req_0 : boolean;
  signal array_obj_ref_2405_index_offset_req_0 : boolean;
  signal array_obj_ref_2405_index_offset_ack_0 : boolean;
  signal array_obj_ref_2405_index_offset_req_1 : boolean;
  signal array_obj_ref_2405_index_offset_ack_1 : boolean;
  signal type_cast_3366_inst_ack_0 : boolean;
  signal addr_of_2406_final_reg_req_0 : boolean;
  signal addr_of_2406_final_reg_ack_0 : boolean;
  signal addr_of_2406_final_reg_req_1 : boolean;
  signal addr_of_2406_final_reg_ack_1 : boolean;
  signal type_cast_3498_inst_req_0 : boolean;
  signal addr_of_3316_final_reg_req_0 : boolean;
  signal type_cast_3327_inst_req_0 : boolean;
  signal addr_of_3316_final_reg_ack_0 : boolean;
  signal ptr_deref_2409_store_0_req_0 : boolean;
  signal ptr_deref_2409_store_0_ack_0 : boolean;
  signal ptr_deref_2409_store_0_req_1 : boolean;
  signal ptr_deref_2409_store_0_ack_1 : boolean;
  signal addr_of_3316_final_reg_req_1 : boolean;
  signal type_cast_2418_inst_req_0 : boolean;
  signal type_cast_2418_inst_ack_0 : boolean;
  signal type_cast_2418_inst_req_1 : boolean;
  signal type_cast_2418_inst_ack_1 : boolean;
  signal addr_of_3316_final_reg_ack_1 : boolean;
  signal type_cast_2482_inst_req_0 : boolean;
  signal type_cast_2482_inst_ack_0 : boolean;
  signal type_cast_2482_inst_req_1 : boolean;
  signal type_cast_2482_inst_ack_1 : boolean;
  signal array_obj_ref_2488_index_offset_req_0 : boolean;
  signal array_obj_ref_2488_index_offset_ack_0 : boolean;
  signal array_obj_ref_2488_index_offset_req_1 : boolean;
  signal array_obj_ref_2488_index_offset_ack_1 : boolean;
  signal addr_of_2489_final_reg_req_0 : boolean;
  signal addr_of_2489_final_reg_ack_0 : boolean;
  signal type_cast_3366_inst_req_1 : boolean;
  signal addr_of_2489_final_reg_req_1 : boolean;
  signal type_cast_3327_inst_ack_0 : boolean;
  signal addr_of_2489_final_reg_ack_1 : boolean;
  signal type_cast_3498_inst_ack_0 : boolean;
  signal type_cast_3327_inst_req_1 : boolean;
  signal type_cast_3327_inst_ack_1 : boolean;
  signal LOAD_pad_3441_load_0_req_0 : boolean;
  signal ptr_deref_2493_load_0_req_0 : boolean;
  signal ptr_deref_2493_load_0_ack_0 : boolean;
  signal LOAD_pad_3441_load_0_ack_0 : boolean;
  signal ptr_deref_2493_load_0_req_1 : boolean;
  signal ptr_deref_2493_load_0_ack_1 : boolean;
  signal type_cast_3309_inst_req_0 : boolean;
  signal type_cast_2507_inst_req_0 : boolean;
  signal type_cast_2507_inst_ack_0 : boolean;
  signal type_cast_3309_inst_ack_0 : boolean;
  signal type_cast_2507_inst_req_1 : boolean;
  signal type_cast_2507_inst_ack_1 : boolean;
  signal type_cast_3498_inst_req_1 : boolean;
  signal type_cast_3366_inst_ack_1 : boolean;
  signal array_obj_ref_2513_index_offset_req_0 : boolean;
  signal array_obj_ref_2513_index_offset_ack_0 : boolean;
  signal array_obj_ref_2513_index_offset_req_1 : boolean;
  signal array_obj_ref_2513_index_offset_ack_1 : boolean;
  signal addr_of_2514_final_reg_req_0 : boolean;
  signal addr_of_2514_final_reg_ack_0 : boolean;
  signal if_stmt_3525_branch_req_0 : boolean;
  signal addr_of_2514_final_reg_req_1 : boolean;
  signal addr_of_2514_final_reg_ack_1 : boolean;
  signal if_stmt_3525_branch_ack_0 : boolean;
  signal type_cast_3309_inst_req_1 : boolean;
  signal type_cast_3498_inst_ack_1 : boolean;
  signal if_stmt_3342_branch_req_0 : boolean;
  signal LOAD_pad_3441_load_0_req_1 : boolean;
  signal ptr_deref_2517_store_0_req_0 : boolean;
  signal ptr_deref_2517_store_0_ack_0 : boolean;
  signal ptr_deref_2517_store_0_req_1 : boolean;
  signal ptr_deref_2517_store_0_ack_1 : boolean;
  signal type_cast_2525_inst_req_0 : boolean;
  signal type_cast_2525_inst_ack_0 : boolean;
  signal type_cast_2525_inst_req_1 : boolean;
  signal type_cast_2525_inst_ack_1 : boolean;
  signal if_stmt_2540_branch_req_0 : boolean;
  signal if_stmt_2540_branch_ack_1 : boolean;
  signal if_stmt_2540_branch_ack_0 : boolean;
  signal type_cast_2564_inst_req_0 : boolean;
  signal type_cast_2564_inst_ack_0 : boolean;
  signal type_cast_2564_inst_req_1 : boolean;
  signal type_cast_2564_inst_ack_1 : boolean;
  signal type_cast_2573_inst_req_0 : boolean;
  signal type_cast_2573_inst_ack_0 : boolean;
  signal type_cast_2573_inst_req_1 : boolean;
  signal type_cast_2573_inst_ack_1 : boolean;
  signal type_cast_2590_inst_req_0 : boolean;
  signal type_cast_2590_inst_ack_0 : boolean;
  signal type_cast_2590_inst_req_1 : boolean;
  signal type_cast_2590_inst_ack_1 : boolean;
  signal if_stmt_2597_branch_req_0 : boolean;
  signal if_stmt_2597_branch_ack_1 : boolean;
  signal if_stmt_2597_branch_ack_0 : boolean;
  signal LOAD_pad_2627_load_0_req_0 : boolean;
  signal LOAD_pad_2627_load_0_ack_0 : boolean;
  signal LOAD_pad_2627_load_0_req_1 : boolean;
  signal LOAD_pad_2627_load_0_ack_1 : boolean;
  signal type_cast_2631_inst_req_0 : boolean;
  signal type_cast_2631_inst_ack_0 : boolean;
  signal type_cast_2631_inst_req_1 : boolean;
  signal type_cast_2631_inst_ack_1 : boolean;
  signal type_cast_2684_inst_req_0 : boolean;
  signal type_cast_2684_inst_ack_0 : boolean;
  signal type_cast_2684_inst_req_1 : boolean;
  signal type_cast_2684_inst_ack_1 : boolean;
  signal if_stmt_2711_branch_req_0 : boolean;
  signal if_stmt_2711_branch_ack_1 : boolean;
  signal if_stmt_2711_branch_ack_0 : boolean;
  signal type_cast_2721_inst_req_0 : boolean;
  signal type_cast_2721_inst_ack_0 : boolean;
  signal type_cast_2721_inst_req_1 : boolean;
  signal type_cast_2721_inst_ack_1 : boolean;
  signal if_stmt_2748_branch_req_0 : boolean;
  signal if_stmt_2748_branch_ack_1 : boolean;
  signal if_stmt_2748_branch_ack_0 : boolean;
  signal type_cast_2758_inst_req_0 : boolean;
  signal type_cast_2758_inst_ack_0 : boolean;
  signal type_cast_2758_inst_req_1 : boolean;
  signal type_cast_2758_inst_ack_1 : boolean;
  signal array_obj_ref_2886_index_offset_req_0 : boolean;
  signal array_obj_ref_2886_index_offset_ack_0 : boolean;
  signal array_obj_ref_2886_index_offset_req_1 : boolean;
  signal array_obj_ref_2886_index_offset_ack_1 : boolean;
  signal addr_of_2887_final_reg_req_0 : boolean;
  signal addr_of_2887_final_reg_ack_0 : boolean;
  signal addr_of_2887_final_reg_req_1 : boolean;
  signal addr_of_2887_final_reg_ack_1 : boolean;
  signal ptr_deref_2891_load_0_req_0 : boolean;
  signal ptr_deref_2891_load_0_ack_0 : boolean;
  signal ptr_deref_2891_load_0_req_1 : boolean;
  signal ptr_deref_2891_load_0_ack_1 : boolean;
  signal type_cast_2905_inst_req_0 : boolean;
  signal type_cast_2905_inst_ack_0 : boolean;
  signal type_cast_2905_inst_req_1 : boolean;
  signal type_cast_2905_inst_ack_1 : boolean;
  signal array_obj_ref_2911_index_offset_req_0 : boolean;
  signal array_obj_ref_2911_index_offset_ack_0 : boolean;
  signal array_obj_ref_2911_index_offset_req_1 : boolean;
  signal array_obj_ref_2911_index_offset_ack_1 : boolean;
  signal addr_of_2912_final_reg_req_0 : boolean;
  signal addr_of_2912_final_reg_ack_0 : boolean;
  signal addr_of_2912_final_reg_req_1 : boolean;
  signal addr_of_2912_final_reg_ack_1 : boolean;
  signal ptr_deref_2915_store_0_req_0 : boolean;
  signal ptr_deref_2915_store_0_ack_0 : boolean;
  signal ptr_deref_2915_store_0_req_1 : boolean;
  signal ptr_deref_2915_store_0_ack_1 : boolean;
  signal type_cast_2923_inst_req_0 : boolean;
  signal type_cast_2923_inst_ack_0 : boolean;
  signal type_cast_2923_inst_req_1 : boolean;
  signal type_cast_2923_inst_ack_1 : boolean;
  signal if_stmt_2938_branch_req_0 : boolean;
  signal if_stmt_2938_branch_ack_1 : boolean;
  signal if_stmt_2938_branch_ack_0 : boolean;
  signal type_cast_2962_inst_req_0 : boolean;
  signal type_cast_2962_inst_ack_0 : boolean;
  signal type_cast_2962_inst_req_1 : boolean;
  signal type_cast_2962_inst_ack_1 : boolean;
  signal type_cast_2971_inst_req_0 : boolean;
  signal type_cast_2971_inst_ack_0 : boolean;
  signal type_cast_2971_inst_req_1 : boolean;
  signal type_cast_2971_inst_ack_1 : boolean;
  signal type_cast_3611_inst_ack_1 : boolean;
  signal ptr_deref_3319_store_0_ack_1 : boolean;
  signal if_stmt_3399_branch_ack_0 : boolean;
  signal if_stmt_3562_branch_ack_0 : boolean;
  signal type_cast_2987_inst_req_0 : boolean;
  signal type_cast_2987_inst_ack_0 : boolean;
  signal type_cast_2987_inst_req_1 : boolean;
  signal type_cast_2987_inst_ack_1 : boolean;
  signal type_cast_3611_inst_req_1 : boolean;
  signal if_stmt_3399_branch_ack_1 : boolean;
  signal if_stmt_2994_branch_req_0 : boolean;
  signal if_stmt_2994_branch_ack_1 : boolean;
  signal if_stmt_3399_branch_req_0 : boolean;
  signal if_stmt_2994_branch_ack_0 : boolean;
  signal array_obj_ref_3315_index_offset_req_1 : boolean;
  signal LOAD_pad_3030_load_0_req_0 : boolean;
  signal ptr_deref_3319_store_0_req_1 : boolean;
  signal LOAD_pad_3030_load_0_ack_0 : boolean;
  signal LOAD_pad_3030_load_0_req_1 : boolean;
  signal LOAD_pad_3030_load_0_ack_1 : boolean;
  signal if_stmt_3562_branch_ack_1 : boolean;
  signal type_cast_3611_inst_ack_0 : boolean;
  signal type_cast_3611_inst_req_0 : boolean;
  signal type_cast_3034_inst_req_0 : boolean;
  signal type_cast_3034_inst_ack_0 : boolean;
  signal if_stmt_3562_branch_req_0 : boolean;
  signal type_cast_3034_inst_req_1 : boolean;
  signal type_cast_3392_inst_ack_1 : boolean;
  signal type_cast_3034_inst_ack_1 : boolean;
  signal if_stmt_3525_branch_ack_1 : boolean;
  signal type_cast_3088_inst_req_0 : boolean;
  signal type_cast_3392_inst_req_1 : boolean;
  signal type_cast_3088_inst_ack_0 : boolean;
  signal type_cast_3088_inst_req_1 : boolean;
  signal type_cast_3088_inst_ack_1 : boolean;
  signal if_stmt_3115_branch_req_0 : boolean;
  signal if_stmt_3115_branch_ack_1 : boolean;
  signal if_stmt_3115_branch_ack_0 : boolean;
  signal type_cast_3445_inst_ack_1 : boolean;
  signal type_cast_3535_inst_ack_1 : boolean;
  signal type_cast_3125_inst_req_0 : boolean;
  signal type_cast_3125_inst_ack_0 : boolean;
  signal if_stmt_3342_branch_ack_0 : boolean;
  signal type_cast_3535_inst_req_1 : boolean;
  signal type_cast_3125_inst_req_1 : boolean;
  signal type_cast_3392_inst_ack_0 : boolean;
  signal type_cast_3125_inst_ack_1 : boolean;
  signal type_cast_3577_inst_ack_1 : boolean;
  signal type_cast_3577_inst_req_1 : boolean;
  signal type_cast_3392_inst_req_0 : boolean;
  signal if_stmt_3152_branch_req_0 : boolean;
  signal type_cast_3309_inst_ack_1 : boolean;
  signal if_stmt_3152_branch_ack_1 : boolean;
  signal if_stmt_3152_branch_ack_0 : boolean;
  signal type_cast_3572_inst_ack_1 : boolean;
  signal if_stmt_3342_branch_ack_1 : boolean;
  signal type_cast_3445_inst_req_1 : boolean;
  signal type_cast_3162_inst_req_0 : boolean;
  signal type_cast_3162_inst_ack_0 : boolean;
  signal type_cast_3535_inst_ack_0 : boolean;
  signal type_cast_3162_inst_req_1 : boolean;
  signal type_cast_3162_inst_ack_1 : boolean;
  signal ptr_deref_3319_store_0_ack_0 : boolean;
  signal type_cast_3572_inst_req_1 : boolean;
  signal type_cast_3535_inst_req_0 : boolean;
  signal type_cast_3167_inst_req_0 : boolean;
  signal type_cast_3167_inst_ack_0 : boolean;
  signal type_cast_3167_inst_req_1 : boolean;
  signal type_cast_3167_inst_ack_1 : boolean;
  signal type_cast_3577_inst_ack_0 : boolean;
  signal type_cast_3577_inst_req_0 : boolean;
  signal type_cast_3445_inst_ack_0 : boolean;
  signal type_cast_3445_inst_req_0 : boolean;
  signal type_cast_3375_inst_ack_1 : boolean;
  signal type_cast_3201_inst_req_0 : boolean;
  signal type_cast_3375_inst_req_1 : boolean;
  signal type_cast_3201_inst_ack_0 : boolean;
  signal type_cast_3201_inst_req_1 : boolean;
  signal type_cast_3201_inst_ack_1 : boolean;
  signal ptr_deref_3319_store_0_req_0 : boolean;
  signal ptr_deref_3295_load_0_ack_1 : boolean;
  signal ptr_deref_3295_load_0_req_1 : boolean;
  signal array_obj_ref_3207_index_offset_req_0 : boolean;
  signal array_obj_ref_3207_index_offset_ack_0 : boolean;
  signal array_obj_ref_3315_index_offset_ack_0 : boolean;
  signal array_obj_ref_3207_index_offset_req_1 : boolean;
  signal type_cast_3375_inst_ack_0 : boolean;
  signal array_obj_ref_3207_index_offset_ack_1 : boolean;
  signal type_cast_3572_inst_ack_0 : boolean;
  signal type_cast_3375_inst_req_0 : boolean;
  signal array_obj_ref_3315_index_offset_req_0 : boolean;
  signal type_cast_3572_inst_req_0 : boolean;
  signal addr_of_3208_final_reg_req_0 : boolean;
  signal addr_of_3208_final_reg_ack_0 : boolean;
  signal addr_of_3208_final_reg_req_1 : boolean;
  signal addr_of_3208_final_reg_ack_1 : boolean;
  signal LOAD_pad_3441_load_0_ack_1 : boolean;
  signal type_cast_1380_inst_req_0 : boolean;
  signal ptr_deref_3211_store_0_req_0 : boolean;
  signal ptr_deref_3211_store_0_ack_0 : boolean;
  signal type_cast_976_inst_req_1 : boolean;
  signal ptr_deref_3211_store_0_req_1 : boolean;
  signal ptr_deref_3211_store_0_ack_1 : boolean;
  signal type_cast_1380_inst_ack_0 : boolean;
  signal type_cast_3220_inst_req_0 : boolean;
  signal type_cast_3220_inst_ack_0 : boolean;
  signal type_cast_978_inst_req_1 : boolean;
  signal type_cast_3220_inst_req_1 : boolean;
  signal type_cast_3220_inst_ack_1 : boolean;
  signal type_cast_978_inst_ack_1 : boolean;
  signal type_cast_3284_inst_req_0 : boolean;
  signal type_cast_1037_inst_req_0 : boolean;
  signal type_cast_3284_inst_ack_0 : boolean;
  signal type_cast_3284_inst_req_1 : boolean;
  signal type_cast_3284_inst_ack_1 : boolean;
  signal array_obj_ref_3290_index_offset_req_0 : boolean;
  signal array_obj_ref_3290_index_offset_ack_0 : boolean;
  signal array_obj_ref_3290_index_offset_req_1 : boolean;
  signal array_obj_ref_3290_index_offset_ack_1 : boolean;
  signal addr_of_3291_final_reg_req_0 : boolean;
  signal addr_of_3291_final_reg_ack_0 : boolean;
  signal addr_of_3291_final_reg_req_1 : boolean;
  signal addr_of_3291_final_reg_ack_1 : boolean;
  signal ptr_deref_3295_load_0_req_0 : boolean;
  signal ptr_deref_3295_load_0_ack_0 : boolean;
  signal array_obj_ref_3617_index_offset_req_0 : boolean;
  signal array_obj_ref_3617_index_offset_ack_0 : boolean;
  signal array_obj_ref_3617_index_offset_req_1 : boolean;
  signal array_obj_ref_3617_index_offset_ack_1 : boolean;
  signal addr_of_3618_final_reg_req_0 : boolean;
  signal addr_of_3618_final_reg_ack_0 : boolean;
  signal addr_of_3618_final_reg_req_1 : boolean;
  signal addr_of_3618_final_reg_ack_1 : boolean;
  signal ptr_deref_3621_store_0_req_0 : boolean;
  signal ptr_deref_3621_store_0_ack_0 : boolean;
  signal ptr_deref_3621_store_0_req_1 : boolean;
  signal ptr_deref_3621_store_0_ack_1 : boolean;
  signal type_cast_3630_inst_req_0 : boolean;
  signal type_cast_3630_inst_ack_0 : boolean;
  signal type_cast_3630_inst_req_1 : boolean;
  signal type_cast_3630_inst_ack_1 : boolean;
  signal type_cast_3694_inst_req_0 : boolean;
  signal type_cast_3694_inst_ack_0 : boolean;
  signal type_cast_3694_inst_req_1 : boolean;
  signal type_cast_3694_inst_ack_1 : boolean;
  signal phi_stmt_979_ack_0 : boolean;
  signal array_obj_ref_3700_index_offset_req_0 : boolean;
  signal array_obj_ref_3700_index_offset_ack_0 : boolean;
  signal array_obj_ref_3700_index_offset_req_1 : boolean;
  signal array_obj_ref_3700_index_offset_ack_1 : boolean;
  signal phi_stmt_973_ack_0 : boolean;
  signal addr_of_3701_final_reg_req_0 : boolean;
  signal addr_of_3701_final_reg_ack_0 : boolean;
  signal addr_of_3701_final_reg_req_1 : boolean;
  signal addr_of_3701_final_reg_ack_1 : boolean;
  signal phi_stmt_1387_req_1 : boolean;
  signal phi_stmt_967_ack_0 : boolean;
  signal type_cast_970_inst_req_0 : boolean;
  signal ptr_deref_3705_load_0_req_0 : boolean;
  signal ptr_deref_3705_load_0_ack_0 : boolean;
  signal phi_stmt_1047_req_1 : boolean;
  signal ptr_deref_3705_load_0_req_1 : boolean;
  signal ptr_deref_3705_load_0_ack_1 : boolean;
  signal type_cast_1053_inst_ack_1 : boolean;
  signal type_cast_978_inst_ack_0 : boolean;
  signal type_cast_3719_inst_req_0 : boolean;
  signal type_cast_1053_inst_req_1 : boolean;
  signal type_cast_3719_inst_ack_0 : boolean;
  signal type_cast_3719_inst_req_1 : boolean;
  signal type_cast_3719_inst_ack_1 : boolean;
  signal phi_stmt_979_req_0 : boolean;
  signal phi_stmt_1047_ack_0 : boolean;
  signal type_cast_978_inst_req_0 : boolean;
  signal type_cast_982_inst_ack_1 : boolean;
  signal type_cast_982_inst_req_1 : boolean;
  signal type_cast_982_inst_ack_0 : boolean;
  signal array_obj_ref_3725_index_offset_req_0 : boolean;
  signal array_obj_ref_3725_index_offset_ack_0 : boolean;
  signal array_obj_ref_3725_index_offset_req_1 : boolean;
  signal type_cast_1053_inst_ack_0 : boolean;
  signal array_obj_ref_3725_index_offset_ack_1 : boolean;
  signal type_cast_982_inst_req_0 : boolean;
  signal type_cast_1053_inst_req_0 : boolean;
  signal addr_of_3726_final_reg_req_0 : boolean;
  signal addr_of_3726_final_reg_ack_0 : boolean;
  signal addr_of_3726_final_reg_req_1 : boolean;
  signal addr_of_3726_final_reg_ack_1 : boolean;
  signal phi_stmt_1040_ack_0 : boolean;
  signal phi_stmt_1034_ack_0 : boolean;
  signal phi_stmt_1047_req_0 : boolean;
  signal phi_stmt_1040_req_0 : boolean;
  signal phi_stmt_1034_req_1 : boolean;
  signal phi_stmt_979_req_1 : boolean;
  signal ptr_deref_3729_store_0_req_0 : boolean;
  signal ptr_deref_3729_store_0_ack_0 : boolean;
  signal ptr_deref_3729_store_0_req_1 : boolean;
  signal ptr_deref_3729_store_0_ack_1 : boolean;
  signal phi_stmt_1381_req_1 : boolean;
  signal type_cast_1386_inst_ack_1 : boolean;
  signal phi_stmt_967_req_0 : boolean;
  signal phi_stmt_1375_req_1 : boolean;
  signal type_cast_1380_inst_ack_1 : boolean;
  signal type_cast_3737_inst_req_0 : boolean;
  signal type_cast_3737_inst_ack_0 : boolean;
  signal type_cast_1039_inst_ack_1 : boolean;
  signal type_cast_3737_inst_req_1 : boolean;
  signal type_cast_3737_inst_ack_1 : boolean;
  signal type_cast_1386_inst_req_1 : boolean;
  signal type_cast_1039_inst_req_1 : boolean;
  signal if_stmt_3752_branch_req_0 : boolean;
  signal type_cast_1380_inst_req_1 : boolean;
  signal if_stmt_3752_branch_ack_1 : boolean;
  signal phi_stmt_973_req_1 : boolean;
  signal if_stmt_3752_branch_ack_0 : boolean;
  signal type_cast_976_inst_ack_0 : boolean;
  signal type_cast_1039_inst_ack_0 : boolean;
  signal type_cast_976_inst_req_0 : boolean;
  signal type_cast_1039_inst_req_0 : boolean;
  signal type_cast_3776_inst_req_0 : boolean;
  signal type_cast_3776_inst_ack_0 : boolean;
  signal type_cast_3776_inst_req_1 : boolean;
  signal type_cast_3776_inst_ack_1 : boolean;
  signal type_cast_1386_inst_ack_0 : boolean;
  signal type_cast_1386_inst_req_0 : boolean;
  signal phi_stmt_1040_req_1 : boolean;
  signal type_cast_3785_inst_req_0 : boolean;
  signal type_cast_1046_inst_ack_1 : boolean;
  signal type_cast_3785_inst_ack_0 : boolean;
  signal type_cast_3785_inst_req_1 : boolean;
  signal type_cast_1046_inst_req_1 : boolean;
  signal type_cast_3785_inst_ack_1 : boolean;
  signal phi_stmt_1034_req_0 : boolean;
  signal type_cast_1037_inst_ack_1 : boolean;
  signal type_cast_3801_inst_req_0 : boolean;
  signal type_cast_3801_inst_ack_0 : boolean;
  signal type_cast_3801_inst_req_1 : boolean;
  signal type_cast_1046_inst_ack_0 : boolean;
  signal type_cast_3801_inst_ack_1 : boolean;
  signal type_cast_1037_inst_req_1 : boolean;
  signal type_cast_970_inst_ack_1 : boolean;
  signal type_cast_970_inst_req_1 : boolean;
  signal if_stmt_3808_branch_req_0 : boolean;
  signal if_stmt_3808_branch_ack_1 : boolean;
  signal if_stmt_3808_branch_ack_0 : boolean;
  signal type_cast_1046_inst_req_0 : boolean;
  signal type_cast_3840_inst_req_0 : boolean;
  signal type_cast_3840_inst_ack_0 : boolean;
  signal type_cast_3840_inst_req_1 : boolean;
  signal type_cast_3840_inst_ack_1 : boolean;
  signal phi_stmt_973_req_0 : boolean;
  signal type_cast_976_inst_ack_1 : boolean;
  signal type_cast_3844_inst_req_0 : boolean;
  signal type_cast_3844_inst_ack_0 : boolean;
  signal type_cast_3844_inst_req_1 : boolean;
  signal type_cast_3844_inst_ack_1 : boolean;
  signal type_cast_970_inst_ack_0 : boolean;
  signal type_cast_1037_inst_ack_0 : boolean;
  signal call_stmt_3857_call_req_0 : boolean;
  signal call_stmt_3857_call_ack_0 : boolean;
  signal call_stmt_3857_call_req_1 : boolean;
  signal call_stmt_3857_call_ack_1 : boolean;
  signal type_cast_3074_inst_ack_0 : boolean;
  signal type_cast_3080_inst_req_1 : boolean;
  signal phi_stmt_3001_req_1 : boolean;
  signal type_cast_3080_inst_req_0 : boolean;
  signal type_cast_3080_inst_ack_0 : boolean;
  signal phi_stmt_338_req_0 : boolean;
  signal type_cast_344_inst_req_0 : boolean;
  signal type_cast_344_inst_ack_0 : boolean;
  signal type_cast_344_inst_req_1 : boolean;
  signal type_cast_344_inst_ack_1 : boolean;
  signal phi_stmt_338_req_1 : boolean;
  signal phi_stmt_338_ack_0 : boolean;
  signal phi_stmt_622_req_0 : boolean;
  signal phi_stmt_630_req_0 : boolean;
  signal phi_stmt_637_req_0 : boolean;
  signal type_cast_629_inst_req_0 : boolean;
  signal type_cast_629_inst_ack_0 : boolean;
  signal type_cast_629_inst_req_1 : boolean;
  signal type_cast_629_inst_ack_1 : boolean;
  signal phi_stmt_622_req_1 : boolean;
  signal type_cast_636_inst_req_0 : boolean;
  signal type_cast_636_inst_ack_0 : boolean;
  signal type_cast_636_inst_req_1 : boolean;
  signal type_cast_636_inst_ack_1 : boolean;
  signal phi_stmt_630_req_1 : boolean;
  signal type_cast_3011_inst_req_0 : boolean;
  signal type_cast_643_inst_req_0 : boolean;
  signal type_cast_643_inst_ack_0 : boolean;
  signal type_cast_643_inst_req_1 : boolean;
  signal type_cast_643_inst_ack_1 : boolean;
  signal phi_stmt_637_req_1 : boolean;
  signal phi_stmt_622_ack_0 : boolean;
  signal phi_stmt_630_ack_0 : boolean;
  signal phi_stmt_637_ack_0 : boolean;
  signal type_cast_972_inst_req_0 : boolean;
  signal type_cast_972_inst_ack_0 : boolean;
  signal type_cast_972_inst_req_1 : boolean;
  signal type_cast_972_inst_ack_1 : boolean;
  signal phi_stmt_967_req_1 : boolean;
  signal type_cast_1378_inst_req_0 : boolean;
  signal type_cast_1378_inst_ack_0 : boolean;
  signal type_cast_1378_inst_req_1 : boolean;
  signal type_cast_1378_inst_ack_1 : boolean;
  signal phi_stmt_1375_req_0 : boolean;
  signal type_cast_1384_inst_req_0 : boolean;
  signal type_cast_1384_inst_ack_0 : boolean;
  signal type_cast_1384_inst_req_1 : boolean;
  signal type_cast_1384_inst_ack_1 : boolean;
  signal phi_stmt_1381_req_0 : boolean;
  signal type_cast_1390_inst_req_0 : boolean;
  signal type_cast_1390_inst_ack_0 : boolean;
  signal type_cast_1390_inst_req_1 : boolean;
  signal type_cast_1390_inst_ack_1 : boolean;
  signal phi_stmt_1387_req_0 : boolean;
  signal phi_stmt_1375_ack_0 : boolean;
  signal phi_stmt_1381_ack_0 : boolean;
  signal phi_stmt_1387_ack_0 : boolean;
  signal type_cast_1454_inst_req_0 : boolean;
  signal type_cast_1454_inst_ack_0 : boolean;
  signal type_cast_1454_inst_req_1 : boolean;
  signal type_cast_1454_inst_ack_1 : boolean;
  signal phi_stmt_1448_req_1 : boolean;
  signal type_cast_1460_inst_req_0 : boolean;
  signal type_cast_1460_inst_ack_0 : boolean;
  signal type_cast_1460_inst_req_1 : boolean;
  signal type_cast_1460_inst_ack_1 : boolean;
  signal phi_stmt_1455_req_1 : boolean;
  signal type_cast_1467_inst_req_0 : boolean;
  signal type_cast_1467_inst_ack_0 : boolean;
  signal type_cast_1467_inst_req_1 : boolean;
  signal type_cast_1467_inst_ack_1 : boolean;
  signal phi_stmt_1461_req_1 : boolean;
  signal phi_stmt_1448_req_0 : boolean;
  signal type_cast_1458_inst_req_0 : boolean;
  signal type_cast_1458_inst_ack_0 : boolean;
  signal type_cast_1458_inst_req_1 : boolean;
  signal type_cast_1458_inst_ack_1 : boolean;
  signal phi_stmt_1455_req_0 : boolean;
  signal phi_stmt_1461_req_0 : boolean;
  signal phi_stmt_1448_ack_0 : boolean;
  signal phi_stmt_1455_ack_0 : boolean;
  signal phi_stmt_1461_ack_0 : boolean;
  signal type_cast_1808_inst_req_0 : boolean;
  signal type_cast_1808_inst_ack_0 : boolean;
  signal type_cast_1808_inst_req_1 : boolean;
  signal type_cast_1808_inst_ack_1 : boolean;
  signal phi_stmt_1803_req_1 : boolean;
  signal type_cast_1802_inst_req_0 : boolean;
  signal type_cast_1802_inst_ack_0 : boolean;
  signal type_cast_1802_inst_req_1 : boolean;
  signal type_cast_1802_inst_ack_1 : boolean;
  signal phi_stmt_1797_req_1 : boolean;
  signal phi_stmt_1790_req_1 : boolean;
  signal type_cast_1806_inst_req_0 : boolean;
  signal type_cast_1806_inst_ack_0 : boolean;
  signal type_cast_1806_inst_req_1 : boolean;
  signal type_cast_1806_inst_ack_1 : boolean;
  signal phi_stmt_1803_req_0 : boolean;
  signal type_cast_1800_inst_req_0 : boolean;
  signal type_cast_1800_inst_ack_0 : boolean;
  signal type_cast_1800_inst_req_1 : boolean;
  signal type_cast_1800_inst_ack_1 : boolean;
  signal phi_stmt_1797_req_0 : boolean;
  signal type_cast_1793_inst_req_0 : boolean;
  signal type_cast_1793_inst_ack_0 : boolean;
  signal type_cast_1793_inst_req_1 : boolean;
  signal type_cast_1793_inst_ack_1 : boolean;
  signal phi_stmt_1790_req_0 : boolean;
  signal phi_stmt_1790_ack_0 : boolean;
  signal phi_stmt_1797_ack_0 : boolean;
  signal phi_stmt_1803_ack_0 : boolean;
  signal type_cast_1863_inst_req_0 : boolean;
  signal type_cast_1863_inst_ack_0 : boolean;
  signal type_cast_1863_inst_req_1 : boolean;
  signal type_cast_1863_inst_ack_1 : boolean;
  signal phi_stmt_1860_req_0 : boolean;
  signal type_cast_1857_inst_req_0 : boolean;
  signal type_cast_1857_inst_ack_0 : boolean;
  signal type_cast_1857_inst_req_1 : boolean;
  signal type_cast_1857_inst_ack_1 : boolean;
  signal phi_stmt_1854_req_0 : boolean;
  signal type_cast_1850_inst_req_0 : boolean;
  signal type_cast_1850_inst_ack_0 : boolean;
  signal type_cast_1850_inst_req_1 : boolean;
  signal type_cast_1850_inst_ack_1 : boolean;
  signal phi_stmt_1847_req_0 : boolean;
  signal type_cast_1865_inst_req_0 : boolean;
  signal type_cast_1865_inst_ack_0 : boolean;
  signal type_cast_1865_inst_req_1 : boolean;
  signal type_cast_1865_inst_ack_1 : boolean;
  signal phi_stmt_1860_req_1 : boolean;
  signal type_cast_1859_inst_req_0 : boolean;
  signal type_cast_1859_inst_ack_0 : boolean;
  signal phi_stmt_3014_ack_0 : boolean;
  signal type_cast_1859_inst_req_1 : boolean;
  signal type_cast_1859_inst_ack_1 : boolean;
  signal phi_stmt_1854_req_1 : boolean;
  signal phi_stmt_3008_ack_0 : boolean;
  signal phi_stmt_1847_req_1 : boolean;
  signal phi_stmt_3001_ack_0 : boolean;
  signal phi_stmt_1847_ack_0 : boolean;
  signal phi_stmt_1854_ack_0 : boolean;
  signal phi_stmt_1860_ack_0 : boolean;
  signal phi_stmt_3008_req_0 : boolean;
  signal type_cast_3074_inst_req_0 : boolean;
  signal phi_stmt_3001_req_0 : boolean;
  signal type_cast_3011_inst_ack_1 : boolean;
  signal type_cast_3004_inst_ack_1 : boolean;
  signal type_cast_3004_inst_req_1 : boolean;
  signal phi_stmt_3071_req_0 : boolean;
  signal type_cast_3011_inst_req_1 : boolean;
  signal type_cast_3004_inst_ack_0 : boolean;
  signal type_cast_3004_inst_req_0 : boolean;
  signal phi_stmt_3077_req_0 : boolean;
  signal type_cast_3074_inst_ack_1 : boolean;
  signal phi_stmt_2187_req_0 : boolean;
  signal type_cast_2199_inst_req_0 : boolean;
  signal type_cast_2199_inst_ack_0 : boolean;
  signal type_cast_2199_inst_req_1 : boolean;
  signal type_cast_2199_inst_ack_1 : boolean;
  signal phi_stmt_2194_req_1 : boolean;
  signal phi_stmt_3014_req_0 : boolean;
  signal type_cast_2203_inst_req_0 : boolean;
  signal type_cast_3017_inst_ack_1 : boolean;
  signal type_cast_2203_inst_ack_0 : boolean;
  signal type_cast_2203_inst_req_1 : boolean;
  signal type_cast_2203_inst_ack_1 : boolean;
  signal phi_stmt_2200_req_0 : boolean;
  signal type_cast_3017_inst_req_1 : boolean;
  signal type_cast_2193_inst_req_0 : boolean;
  signal type_cast_2193_inst_ack_0 : boolean;
  signal type_cast_2193_inst_req_1 : boolean;
  signal type_cast_2193_inst_ack_1 : boolean;
  signal phi_stmt_2187_req_1 : boolean;
  signal type_cast_3017_inst_ack_0 : boolean;
  signal type_cast_2197_inst_req_0 : boolean;
  signal type_cast_2197_inst_ack_0 : boolean;
  signal type_cast_3017_inst_req_0 : boolean;
  signal type_cast_2197_inst_req_1 : boolean;
  signal type_cast_2197_inst_ack_1 : boolean;
  signal phi_stmt_2194_req_0 : boolean;
  signal phi_stmt_3064_req_1 : boolean;
  signal type_cast_2205_inst_req_0 : boolean;
  signal type_cast_2205_inst_ack_0 : boolean;
  signal type_cast_2205_inst_req_1 : boolean;
  signal type_cast_2205_inst_ack_1 : boolean;
  signal phi_stmt_2200_req_1 : boolean;
  signal phi_stmt_3008_req_1 : boolean;
  signal type_cast_3013_inst_ack_1 : boolean;
  signal type_cast_3070_inst_ack_1 : boolean;
  signal type_cast_3074_inst_req_1 : boolean;
  signal phi_stmt_2187_ack_0 : boolean;
  signal phi_stmt_2194_ack_0 : boolean;
  signal phi_stmt_2200_ack_0 : boolean;
  signal type_cast_3011_inst_ack_0 : boolean;
  signal type_cast_3013_inst_req_1 : boolean;
  signal type_cast_3080_inst_ack_1 : boolean;
  signal type_cast_3070_inst_req_1 : boolean;
  signal type_cast_2268_inst_req_0 : boolean;
  signal type_cast_2268_inst_ack_0 : boolean;
  signal phi_stmt_3014_req_1 : boolean;
  signal type_cast_2268_inst_req_1 : boolean;
  signal type_cast_3019_inst_ack_1 : boolean;
  signal type_cast_2268_inst_ack_1 : boolean;
  signal phi_stmt_2262_req_1 : boolean;
  signal type_cast_3013_inst_ack_0 : boolean;
  signal type_cast_3070_inst_ack_0 : boolean;
  signal type_cast_3070_inst_req_0 : boolean;
  signal type_cast_2274_inst_req_0 : boolean;
  signal type_cast_2274_inst_ack_0 : boolean;
  signal type_cast_3019_inst_req_1 : boolean;
  signal type_cast_2274_inst_req_1 : boolean;
  signal type_cast_2274_inst_ack_1 : boolean;
  signal phi_stmt_2269_req_1 : boolean;
  signal type_cast_3013_inst_req_0 : boolean;
  signal type_cast_2281_inst_req_0 : boolean;
  signal type_cast_2281_inst_ack_0 : boolean;
  signal type_cast_2281_inst_req_1 : boolean;
  signal type_cast_3019_inst_ack_0 : boolean;
  signal type_cast_2281_inst_ack_1 : boolean;
  signal phi_stmt_2275_req_1 : boolean;
  signal type_cast_3019_inst_req_0 : boolean;
  signal phi_stmt_2262_req_0 : boolean;
  signal type_cast_2272_inst_req_0 : boolean;
  signal type_cast_2272_inst_ack_0 : boolean;
  signal type_cast_2272_inst_req_1 : boolean;
  signal type_cast_2272_inst_ack_1 : boolean;
  signal phi_stmt_2269_req_0 : boolean;
  signal phi_stmt_2275_req_0 : boolean;
  signal phi_stmt_2262_ack_0 : boolean;
  signal phi_stmt_2269_ack_0 : boolean;
  signal phi_stmt_2275_ack_0 : boolean;
  signal phi_stmt_2604_req_1 : boolean;
  signal type_cast_2616_inst_req_0 : boolean;
  signal type_cast_2616_inst_ack_0 : boolean;
  signal type_cast_2616_inst_req_1 : boolean;
  signal type_cast_2616_inst_ack_1 : boolean;
  signal phi_stmt_2611_req_1 : boolean;
  signal type_cast_2622_inst_req_0 : boolean;
  signal type_cast_2622_inst_ack_0 : boolean;
  signal type_cast_2622_inst_req_1 : boolean;
  signal type_cast_2622_inst_ack_1 : boolean;
  signal phi_stmt_2617_req_1 : boolean;
  signal type_cast_2607_inst_req_0 : boolean;
  signal type_cast_2607_inst_ack_0 : boolean;
  signal type_cast_2607_inst_req_1 : boolean;
  signal type_cast_2607_inst_ack_1 : boolean;
  signal phi_stmt_2604_req_0 : boolean;
  signal type_cast_2614_inst_req_0 : boolean;
  signal type_cast_2614_inst_ack_0 : boolean;
  signal type_cast_2614_inst_req_1 : boolean;
  signal type_cast_2614_inst_ack_1 : boolean;
  signal phi_stmt_2611_req_0 : boolean;
  signal type_cast_2620_inst_req_0 : boolean;
  signal type_cast_2620_inst_ack_0 : boolean;
  signal type_cast_2620_inst_req_1 : boolean;
  signal type_cast_2620_inst_ack_1 : boolean;
  signal phi_stmt_2617_req_0 : boolean;
  signal phi_stmt_2604_ack_0 : boolean;
  signal phi_stmt_2611_ack_0 : boolean;
  signal phi_stmt_2617_ack_0 : boolean;
  signal type_cast_2667_inst_req_0 : boolean;
  signal type_cast_2667_inst_ack_0 : boolean;
  signal type_cast_2667_inst_req_1 : boolean;
  signal type_cast_2667_inst_ack_1 : boolean;
  signal phi_stmt_2661_req_1 : boolean;
  signal type_cast_2673_inst_req_0 : boolean;
  signal type_cast_2673_inst_ack_0 : boolean;
  signal type_cast_2673_inst_req_1 : boolean;
  signal type_cast_2673_inst_ack_1 : boolean;
  signal phi_stmt_2668_req_1 : boolean;
  signal type_cast_2679_inst_req_0 : boolean;
  signal type_cast_2679_inst_ack_0 : boolean;
  signal type_cast_2679_inst_req_1 : boolean;
  signal type_cast_2679_inst_ack_1 : boolean;
  signal phi_stmt_2674_req_1 : boolean;
  signal phi_stmt_2661_req_0 : boolean;
  signal type_cast_2671_inst_req_0 : boolean;
  signal type_cast_2671_inst_ack_0 : boolean;
  signal type_cast_2671_inst_req_1 : boolean;
  signal type_cast_2671_inst_ack_1 : boolean;
  signal phi_stmt_2668_req_0 : boolean;
  signal type_cast_2677_inst_req_0 : boolean;
  signal type_cast_2677_inst_ack_0 : boolean;
  signal type_cast_2677_inst_req_1 : boolean;
  signal type_cast_2677_inst_ack_1 : boolean;
  signal phi_stmt_2674_req_0 : boolean;
  signal phi_stmt_2661_ack_0 : boolean;
  signal phi_stmt_2668_ack_0 : boolean;
  signal phi_stmt_2674_ack_0 : boolean;
  signal phi_stmt_3077_req_1 : boolean;
  signal phi_stmt_3064_req_0 : boolean;
  signal type_cast_3076_inst_req_0 : boolean;
  signal type_cast_3076_inst_ack_0 : boolean;
  signal type_cast_3076_inst_req_1 : boolean;
  signal type_cast_3076_inst_ack_1 : boolean;
  signal phi_stmt_3071_req_1 : boolean;
  signal phi_stmt_3064_ack_0 : boolean;
  signal phi_stmt_3071_ack_0 : boolean;
  signal phi_stmt_3077_ack_0 : boolean;
  signal type_cast_3422_inst_req_0 : boolean;
  signal type_cast_3422_inst_ack_0 : boolean;
  signal type_cast_3422_inst_req_1 : boolean;
  signal type_cast_3422_inst_ack_1 : boolean;
  signal phi_stmt_3419_req_0 : boolean;
  signal phi_stmt_3406_req_0 : boolean;
  signal type_cast_3416_inst_req_0 : boolean;
  signal type_cast_3416_inst_ack_0 : boolean;
  signal type_cast_3416_inst_req_1 : boolean;
  signal type_cast_3416_inst_ack_1 : boolean;
  signal phi_stmt_3413_req_0 : boolean;
  signal type_cast_3424_inst_req_0 : boolean;
  signal type_cast_3424_inst_ack_0 : boolean;
  signal type_cast_3424_inst_req_1 : boolean;
  signal type_cast_3424_inst_ack_1 : boolean;
  signal phi_stmt_3419_req_1 : boolean;
  signal type_cast_3412_inst_req_0 : boolean;
  signal type_cast_3412_inst_ack_0 : boolean;
  signal type_cast_3412_inst_req_1 : boolean;
  signal type_cast_3412_inst_ack_1 : boolean;
  signal phi_stmt_3406_req_1 : boolean;
  signal type_cast_3418_inst_req_0 : boolean;
  signal type_cast_3418_inst_ack_0 : boolean;
  signal type_cast_3418_inst_req_1 : boolean;
  signal type_cast_3418_inst_ack_1 : boolean;
  signal phi_stmt_3413_req_1 : boolean;
  signal phi_stmt_3406_ack_0 : boolean;
  signal phi_stmt_3413_ack_0 : boolean;
  signal phi_stmt_3419_ack_0 : boolean;
  signal type_cast_3481_inst_req_0 : boolean;
  signal type_cast_3481_inst_ack_0 : boolean;
  signal type_cast_3481_inst_req_1 : boolean;
  signal type_cast_3481_inst_ack_1 : boolean;
  signal phi_stmt_3475_req_1 : boolean;
  signal type_cast_3487_inst_req_0 : boolean;
  signal type_cast_3487_inst_ack_0 : boolean;
  signal type_cast_3487_inst_req_1 : boolean;
  signal type_cast_3487_inst_ack_1 : boolean;
  signal phi_stmt_3482_req_1 : boolean;
  signal type_cast_3493_inst_req_0 : boolean;
  signal type_cast_3493_inst_ack_0 : boolean;
  signal type_cast_3493_inst_req_1 : boolean;
  signal type_cast_3493_inst_ack_1 : boolean;
  signal phi_stmt_3488_req_1 : boolean;
  signal phi_stmt_3475_req_0 : boolean;
  signal type_cast_3485_inst_req_0 : boolean;
  signal type_cast_3485_inst_ack_0 : boolean;
  signal type_cast_3485_inst_req_1 : boolean;
  signal type_cast_3485_inst_ack_1 : boolean;
  signal phi_stmt_3482_req_0 : boolean;
  signal type_cast_3491_inst_req_0 : boolean;
  signal type_cast_3491_inst_ack_0 : boolean;
  signal type_cast_3491_inst_req_1 : boolean;
  signal type_cast_3491_inst_ack_1 : boolean;
  signal phi_stmt_3488_req_0 : boolean;
  signal phi_stmt_3475_ack_0 : boolean;
  signal phi_stmt_3482_ack_0 : boolean;
  signal phi_stmt_3488_ack_0 : boolean;
  signal phi_stmt_3815_req_0 : boolean;
  signal type_cast_3827_inst_req_0 : boolean;
  signal type_cast_3827_inst_ack_0 : boolean;
  signal type_cast_3827_inst_req_1 : boolean;
  signal type_cast_3827_inst_ack_1 : boolean;
  signal phi_stmt_3822_req_1 : boolean;
  signal type_cast_3831_inst_req_0 : boolean;
  signal type_cast_3831_inst_ack_0 : boolean;
  signal type_cast_3831_inst_req_1 : boolean;
  signal type_cast_3831_inst_ack_1 : boolean;
  signal phi_stmt_3828_req_0 : boolean;
  signal type_cast_3821_inst_req_0 : boolean;
  signal type_cast_3821_inst_ack_0 : boolean;
  signal type_cast_3821_inst_req_1 : boolean;
  signal type_cast_3821_inst_ack_1 : boolean;
  signal phi_stmt_3815_req_1 : boolean;
  signal type_cast_3825_inst_req_0 : boolean;
  signal type_cast_3825_inst_ack_0 : boolean;
  signal type_cast_3825_inst_req_1 : boolean;
  signal type_cast_3825_inst_ack_1 : boolean;
  signal phi_stmt_3822_req_0 : boolean;
  signal type_cast_3833_inst_req_0 : boolean;
  signal type_cast_3833_inst_ack_0 : boolean;
  signal type_cast_3833_inst_req_1 : boolean;
  signal type_cast_3833_inst_ack_1 : boolean;
  signal phi_stmt_3828_req_1 : boolean;
  signal phi_stmt_3815_ack_0 : boolean;
  signal phi_stmt_3822_ack_0 : boolean;
  signal phi_stmt_3828_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_CP_676_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_676_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_CP_676_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_676_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_CP_676: Block -- control-path 
    signal zeropad3D_CP_676_elements: BooleanArray(956 downto 0);
    -- 
  begin -- 
    zeropad3D_CP_676_elements(0) <= zeropad3D_CP_676_start;
    zeropad3D_CP_676_symbol <= zeropad3D_CP_676_elements(577);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	31 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	35 
    -- CP-element group 0:  members (24) 
      -- CP-element group 0: 	 branch_block_stmt_223/branch_block_stmt_223__entry__
      -- CP-element group 0: 	 branch_block_stmt_223/$entry
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/$entry
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_update_start_
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_update_start_
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_update_start_
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_update_start_
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_Update/cr
      -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => RPIPE_zeropad_input_pipe_225_inst_req_0); -- 
    cr_1160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => STORE_pad_242_store_0_req_1); -- 
    cr_1216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_256_inst_req_1); -- 
    cr_1230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_260_inst_req_1); -- 
    cr_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_264_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	628 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	589 
    -- CP-element group 1: 	590 
    -- CP-element group 1: 	592 
    -- CP-element group 1: 	593 
    -- CP-element group 1: 	595 
    -- CP-element group 1: 	596 
    -- CP-element group 1:  members (27) 
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_223/merge_stmt_966__exit__
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/SplitProtocol/Update/cr
      -- 
    rr_6755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(1), ack => type_cast_629_inst_req_0); -- 
    cr_6760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(1), ack => type_cast_629_inst_req_1); -- 
    rr_6778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(1), ack => type_cast_636_inst_req_0); -- 
    cr_6783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(1), ack => type_cast_636_inst_req_1); -- 
    rr_6801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(1), ack => type_cast_643_inst_req_0); -- 
    cr_6806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(1), ack => type_cast_643_inst_req_1); -- 
    zeropad3D_CP_676_elements(1) <= zeropad3D_CP_676_elements(628);
    -- CP-element group 2:  merge  fork  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	674 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	629 
    -- CP-element group 2: 	630 
    -- CP-element group 2: 	632 
    -- CP-element group 2: 	633 
    -- CP-element group 2: 	635 
    -- CP-element group 2: 	636 
    -- CP-element group 2:  members (27) 
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313
      -- CP-element group 2: 	 branch_block_stmt_223/merge_stmt_1374__exit__
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/SplitProtocol/$entry
      -- 
    cr_7099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(2), ack => type_cast_1053_inst_req_1); -- 
    rr_7094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(2), ack => type_cast_1053_inst_req_0); -- 
    cr_7053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(2), ack => type_cast_1039_inst_req_1); -- 
    rr_7048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(2), ack => type_cast_1039_inst_req_0); -- 
    cr_7076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(2), ack => type_cast_1046_inst_req_1); -- 
    rr_7071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(2), ack => type_cast_1046_inst_req_0); -- 
    zeropad3D_CP_676_elements(2) <= zeropad3D_CP_676_elements(674);
    -- CP-element group 3:  merge  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	720 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	675 
    -- CP-element group 3: 	676 
    -- CP-element group 3: 	678 
    -- CP-element group 3: 	679 
    -- CP-element group 3: 	681 
    -- CP-element group 3: 	682 
    -- CP-element group 3:  members (27) 
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529
      -- CP-element group 3: 	 branch_block_stmt_223/merge_stmt_1789__exit__
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/SplitProtocol/Update/cr
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/SplitProtocol/Update/cr
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Update/cr
      -- 
    rr_7383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(3), ack => type_cast_1454_inst_req_0); -- 
    cr_7388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(3), ack => type_cast_1454_inst_req_1); -- 
    rr_7406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(3), ack => type_cast_1460_inst_req_0); -- 
    cr_7411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(3), ack => type_cast_1460_inst_req_1); -- 
    rr_7429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(3), ack => type_cast_1467_inst_req_0); -- 
    cr_7434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(3), ack => type_cast_1467_inst_req_1); -- 
    zeropad3D_CP_676_elements(3) <= zeropad3D_CP_676_elements(720);
    -- CP-element group 4:  merge  fork  transition  place  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	768 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	721 
    -- CP-element group 4: 	722 
    -- CP-element group 4: 	724 
    -- CP-element group 4: 	725 
    -- CP-element group 4: 	727 
    -- CP-element group 4: 	728 
    -- CP-element group 4:  members (27) 
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751
      -- CP-element group 4: 	 branch_block_stmt_223/merge_stmt_2186__exit__
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/SplitProtocol/Update/cr
      -- 
    rr_7718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(4), ack => type_cast_1863_inst_req_0); -- 
    cr_7723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(4), ack => type_cast_1863_inst_req_1); -- 
    rr_7741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(4), ack => type_cast_1857_inst_req_0); -- 
    cr_7746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(4), ack => type_cast_1857_inst_req_1); -- 
    rr_7764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(4), ack => type_cast_1850_inst_req_0); -- 
    cr_7769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(4), ack => type_cast_1850_inst_req_1); -- 
    zeropad3D_CP_676_elements(4) <= zeropad3D_CP_676_elements(768);
    -- CP-element group 5:  merge  fork  transition  place  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	814 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	769 
    -- CP-element group 5: 	770 
    -- CP-element group 5: 	772 
    -- CP-element group 5: 	773 
    -- CP-element group 5: 	775 
    -- CP-element group 5: 	776 
    -- CP-element group 5:  members (27) 
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967
      -- CP-element group 5: 	 branch_block_stmt_223/merge_stmt_2603__exit__
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/SplitProtocol/Update/cr
      -- 
    rr_8068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(5), ack => type_cast_2268_inst_req_0); -- 
    cr_8073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(5), ack => type_cast_2268_inst_req_1); -- 
    rr_8091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(5), ack => type_cast_2274_inst_req_0); -- 
    cr_8096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(5), ack => type_cast_2274_inst_req_1); -- 
    rr_8114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(5), ack => type_cast_2281_inst_req_0); -- 
    cr_8119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(5), ack => type_cast_2281_inst_req_1); -- 
    zeropad3D_CP_676_elements(5) <= zeropad3D_CP_676_elements(814);
    -- CP-element group 6:  merge  fork  transition  place  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	862 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	815 
    -- CP-element group 6: 	816 
    -- CP-element group 6: 	818 
    -- CP-element group 6: 	819 
    -- CP-element group 6: 	821 
    -- CP-element group 6: 	822 
    -- CP-element group 6:  members (27) 
      -- CP-element group 6: 	 branch_block_stmt_223/merge_stmt_3000__exit__
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/SplitProtocol/Update/cr
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/SplitProtocol/Update/cr
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/SplitProtocol/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/SplitProtocol/Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/SplitProtocol/Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/SplitProtocol/Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/SplitProtocol/Update/cr
      -- 
    rr_8403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => type_cast_2667_inst_req_0); -- 
    cr_8408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => type_cast_2667_inst_req_1); -- 
    rr_8426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => type_cast_2673_inst_req_0); -- 
    cr_8431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => type_cast_2673_inst_req_1); -- 
    rr_8449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => type_cast_2679_inst_req_0); -- 
    cr_8454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => type_cast_2679_inst_req_1); -- 
    zeropad3D_CP_676_elements(6) <= zeropad3D_CP_676_elements(862);
    -- CP-element group 7:  merge  fork  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	908 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	863 
    -- CP-element group 7: 	864 
    -- CP-element group 7: 	866 
    -- CP-element group 7: 	867 
    -- CP-element group 7: 	869 
    -- CP-element group 7: 	870 
    -- CP-element group 7:  members (27) 
      -- CP-element group 7: 	 branch_block_stmt_223/merge_stmt_3405__exit__
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/SplitProtocol/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/$entry
      -- 
    cr_8758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(7), ack => type_cast_3080_inst_req_1); -- 
    rr_8753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(7), ack => type_cast_3080_inst_req_0); -- 
    rr_8799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(7), ack => type_cast_3074_inst_req_0); -- 
    cr_8804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(7), ack => type_cast_3074_inst_req_1); -- 
    cr_8781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(7), ack => type_cast_3070_inst_req_1); -- 
    rr_8776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(7), ack => type_cast_3070_inst_req_0); -- 
    zeropad3D_CP_676_elements(7) <= zeropad3D_CP_676_elements(908);
    -- CP-element group 8:  merge  fork  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	956 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	909 
    -- CP-element group 8: 	910 
    -- CP-element group 8: 	912 
    -- CP-element group 8: 	913 
    -- CP-element group 8: 	915 
    -- CP-element group 8: 	916 
    -- CP-element group 8:  members (27) 
      -- CP-element group 8: 	 branch_block_stmt_223/merge_stmt_3814__exit__
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/SplitProtocol/Update/cr
      -- 
    rr_9088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => type_cast_3481_inst_req_0); -- 
    cr_9093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => type_cast_3481_inst_req_1); -- 
    rr_9111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => type_cast_3487_inst_req_0); -- 
    cr_9116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => type_cast_3487_inst_req_1); -- 
    rr_9134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => type_cast_3493_inst_req_0); -- 
    cr_9139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => type_cast_3493_inst_req_1); -- 
    zeropad3D_CP_676_elements(8) <= zeropad3D_CP_676_elements(956);
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_update_start_
      -- CP-element group 9: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_Update/cr
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_225_inst_ack_0, ack => zeropad3D_CP_676_elements(9)); -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(9), ack => RPIPE_zeropad_input_pipe_225_inst_req_1); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_225_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_Sample/rr
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_225_inst_ack_1, ack => zeropad3D_CP_676_elements(10)); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(10), ack => RPIPE_zeropad_input_pipe_228_inst_req_0); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_update_start_
      -- CP-element group 11: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_Update/cr
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_228_inst_ack_0, ack => zeropad3D_CP_676_elements(11)); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(11), ack => RPIPE_zeropad_input_pipe_228_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_228_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_Sample/rr
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_228_inst_ack_1, ack => zeropad3D_CP_676_elements(12)); -- 
    rr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(12), ack => RPIPE_zeropad_input_pipe_231_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_update_start_
      -- CP-element group 13: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_Update/cr
      -- 
    ra_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_231_inst_ack_0, ack => zeropad3D_CP_676_elements(13)); -- 
    cr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(13), ack => RPIPE_zeropad_input_pipe_231_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	30 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_231_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_Sample/rr
      -- 
    ca_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_231_inst_ack_1, ack => zeropad3D_CP_676_elements(14)); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(14), ack => RPIPE_zeropad_input_pipe_234_inst_req_0); -- 
    rr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(14), ack => type_cast_256_inst_req_0); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_update_start_
      -- CP-element group 15: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_Update/cr
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_234_inst_ack_0, ack => zeropad3D_CP_676_elements(15)); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(15), ack => RPIPE_zeropad_input_pipe_234_inst_req_1); -- 
    -- CP-element group 16:  fork  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16: 	32 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_234_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_Sample/rr
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_234_inst_ack_1, ack => zeropad3D_CP_676_elements(16)); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(16), ack => RPIPE_zeropad_input_pipe_237_inst_req_0); -- 
    rr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(16), ack => type_cast_260_inst_req_0); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_update_start_
      -- CP-element group 17: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_Update/cr
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_237_inst_ack_0, ack => zeropad3D_CP_676_elements(17)); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(17), ack => RPIPE_zeropad_input_pipe_237_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	34 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_237_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_Sample/rr
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_237_inst_ack_1, ack => zeropad3D_CP_676_elements(18)); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(18), ack => RPIPE_zeropad_input_pipe_240_inst_req_0); -- 
    rr_1239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(18), ack => type_cast_264_inst_req_0); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_update_start_
      -- CP-element group 19: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_Update/cr
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_240_inst_ack_0, ack => zeropad3D_CP_676_elements(19)); -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(19), ack => RPIPE_zeropad_input_pipe_240_inst_req_1); -- 
    -- CP-element group 20:  fork  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20: 	24 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_240_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_Sample/rr
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_240_inst_ack_1, ack => zeropad3D_CP_676_elements(20)); -- 
    rr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(20), ack => RPIPE_zeropad_input_pipe_246_inst_req_0); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/STORE_pad_242_Split/$entry
      -- CP-element group 21: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/STORE_pad_242_Split/$exit
      -- CP-element group 21: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/STORE_pad_242_Split/split_req
      -- CP-element group 21: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/STORE_pad_242_Split/split_ack
      -- CP-element group 21: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/word_access_start/$entry
      -- CP-element group 21: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/word_access_start/word_0/$entry
      -- CP-element group 21: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/word_access_start/word_0/rr
      -- 
    rr_1149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(21), ack => STORE_pad_242_store_0_req_0); -- 
    zeropad3D_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(0) & zeropad3D_CP_676_elements(20);
      gj_zeropad3D_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/word_access_start/$exit
      -- CP-element group 22: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/word_access_start/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Sample/word_access_start/word_0/ra
      -- 
    ra_1150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_242_store_0_ack_0, ack => zeropad3D_CP_676_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	36 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Update/word_access_complete/$exit
      -- CP-element group 23: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Update/word_access_complete/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/STORE_pad_242_Update/word_access_complete/word_0/ca
      -- 
    ca_1161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_pad_242_store_0_ack_1, ack => zeropad3D_CP_676_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	20 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_update_start_
      -- CP-element group 24: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_Update/cr
      -- 
    ra_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_246_inst_ack_0, ack => zeropad3D_CP_676_elements(24)); -- 
    cr_1174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(24), ack => RPIPE_zeropad_input_pipe_246_inst_req_1); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_246_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_Sample/rr
      -- 
    ca_1175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_246_inst_ack_1, ack => zeropad3D_CP_676_elements(25)); -- 
    rr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(25), ack => RPIPE_zeropad_input_pipe_249_inst_req_0); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_update_start_
      -- CP-element group 26: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_Update/cr
      -- 
    ra_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_249_inst_ack_0, ack => zeropad3D_CP_676_elements(26)); -- 
    cr_1188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(26), ack => RPIPE_zeropad_input_pipe_249_inst_req_1); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_249_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_Sample/rr
      -- 
    ca_1189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_249_inst_ack_1, ack => zeropad3D_CP_676_elements(27)); -- 
    rr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(27), ack => RPIPE_zeropad_input_pipe_252_inst_req_0); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_update_start_
      -- CP-element group 28: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_Update/cr
      -- 
    ra_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_252_inst_ack_0, ack => zeropad3D_CP_676_elements(28)); -- 
    cr_1202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(28), ack => RPIPE_zeropad_input_pipe_252_inst_req_1); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	36 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/RPIPE_zeropad_input_pipe_252_Update/ca
      -- 
    ca_1203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_252_inst_ack_1, ack => zeropad3D_CP_676_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	14 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_Sample/ra
      -- 
    ra_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_256_inst_ack_0, ack => zeropad3D_CP_676_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	0 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	36 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_256_Update/ca
      -- 
    ca_1217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_256_inst_ack_1, ack => zeropad3D_CP_676_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	16 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_Sample/ra
      -- 
    ra_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_0, ack => zeropad3D_CP_676_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_260_Update/ca
      -- 
    ca_1231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_1, ack => zeropad3D_CP_676_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	18 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_Sample/ra
      -- 
    ra_1240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_264_inst_ack_0, ack => zeropad3D_CP_676_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	0 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/type_cast_264_Update/ca
      -- 
    ca_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_264_inst_ack_1, ack => zeropad3D_CP_676_elements(35)); -- 
    -- CP-element group 36:  branch  join  transition  place  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	23 
    -- CP-element group 36: 	29 
    -- CP-element group 36: 	31 
    -- CP-element group 36: 	33 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (10) 
      -- CP-element group 36: 	 branch_block_stmt_223/if_stmt_288__entry__
      -- CP-element group 36: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287__exit__
      -- CP-element group 36: 	 branch_block_stmt_223/assign_stmt_226_to_assign_stmt_287/$exit
      -- CP-element group 36: 	 branch_block_stmt_223/if_stmt_288_dead_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_223/if_stmt_288_eval_test/$entry
      -- CP-element group 36: 	 branch_block_stmt_223/if_stmt_288_eval_test/$exit
      -- CP-element group 36: 	 branch_block_stmt_223/if_stmt_288_eval_test/branch_req
      -- CP-element group 36: 	 branch_block_stmt_223/R_cmp1840_289_place
      -- CP-element group 36: 	 branch_block_stmt_223/if_stmt_288_if_link/$entry
      -- CP-element group 36: 	 branch_block_stmt_223/if_stmt_288_else_link/$entry
      -- 
    branch_req_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(36), ack => if_stmt_288_branch_req_0); -- 
    zeropad3D_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(23) & zeropad3D_CP_676_elements(29) & zeropad3D_CP_676_elements(31) & zeropad3D_CP_676_elements(33) & zeropad3D_CP_676_elements(35);
      gj_zeropad3D_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  place  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	584 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 branch_block_stmt_223/if_stmt_288_if_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_223/if_stmt_288_if_link/if_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_223/entry_forx_xend
      -- CP-element group 37: 	 branch_block_stmt_223/entry_forx_xend_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_223/entry_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_288_branch_ack_1, ack => zeropad3D_CP_676_elements(37)); -- 
    -- CP-element group 38:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	40 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	42 
    -- CP-element group 38: 	43 
    -- CP-element group 38: 	44 
    -- CP-element group 38:  members (30) 
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335__entry__
      -- CP-element group 38: 	 branch_block_stmt_223/merge_stmt_294__exit__
      -- CP-element group 38: 	 branch_block_stmt_223/if_stmt_288_else_link/$exit
      -- CP-element group 38: 	 branch_block_stmt_223/if_stmt_288_else_link/else_choice_transition
      -- CP-element group 38: 	 branch_block_stmt_223/entry_bbx_xnph
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/$entry
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_update_start_
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_Update/cr
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_update_start_
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_Update/cr
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_update_start_
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_Update/cr
      -- CP-element group 38: 	 branch_block_stmt_223/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_223/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 38: 	 branch_block_stmt_223/merge_stmt_294_PhiReqMerge
      -- CP-element group 38: 	 branch_block_stmt_223/merge_stmt_294_PhiAck/$entry
      -- CP-element group 38: 	 branch_block_stmt_223/merge_stmt_294_PhiAck/$exit
      -- CP-element group 38: 	 branch_block_stmt_223/merge_stmt_294_PhiAck/dummy
      -- 
    else_choice_transition_1262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_288_branch_ack_0, ack => zeropad3D_CP_676_elements(38)); -- 
    rr_1275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(38), ack => type_cast_297_inst_req_0); -- 
    cr_1280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(38), ack => type_cast_297_inst_req_1); -- 
    rr_1289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(38), ack => type_cast_301_inst_req_0); -- 
    cr_1294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(38), ack => type_cast_301_inst_req_1); -- 
    rr_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(38), ack => type_cast_310_inst_req_0); -- 
    cr_1308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(38), ack => type_cast_310_inst_req_1); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_Sample/ra
      -- 
    ra_1276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_297_inst_ack_0, ack => zeropad3D_CP_676_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	45 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_297_Update/ca
      -- 
    ca_1281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_297_inst_ack_1, ack => zeropad3D_CP_676_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_Sample/ra
      -- 
    ra_1290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_301_inst_ack_0, ack => zeropad3D_CP_676_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	38 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_301_Update/ca
      -- 
    ca_1295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_301_inst_ack_1, ack => zeropad3D_CP_676_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	38 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_Sample/ra
      -- 
    ra_1304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_310_inst_ack_0, ack => zeropad3D_CP_676_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	38 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/type_cast_310_Update/ca
      -- 
    ca_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_310_inst_ack_1, ack => zeropad3D_CP_676_elements(44)); -- 
    -- CP-element group 45:  join  transition  place  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	40 
    -- CP-element group 45: 	42 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	578 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_223/bbx_xnph_forx_xbody
      -- CP-element group 45: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335__exit__
      -- CP-element group 45: 	 branch_block_stmt_223/assign_stmt_298_to_assign_stmt_335/$exit
      -- CP-element group 45: 	 branch_block_stmt_223/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 45: 	 branch_block_stmt_223/bbx_xnph_forx_xbody_PhiReq/phi_stmt_338/$entry
      -- CP-element group 45: 	 branch_block_stmt_223/bbx_xnph_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/$entry
      -- 
    zeropad3D_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(40) & zeropad3D_CP_676_elements(42) & zeropad3D_CP_676_elements(44);
      gj_zeropad3D_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	583 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	85 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_final_index_sum_regn_sample_complete
      -- CP-element group 46: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_final_index_sum_regn_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_final_index_sum_regn_Sample/ack
      -- 
    ack_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_350_index_offset_ack_0, ack => zeropad3D_CP_676_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	583 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (11) 
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_root_address_calculated
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_offset_calculated
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_final_index_sum_regn_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_final_index_sum_regn_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_base_plus_offset/$entry
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_base_plus_offset/$exit
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_base_plus_offset/sum_rename_req
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_base_plus_offset/sum_rename_ack
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_request/$entry
      -- CP-element group 47: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_request/req
      -- 
    ack_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_350_index_offset_ack_1, ack => zeropad3D_CP_676_elements(47)); -- 
    req_1352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(47), ack => addr_of_351_final_reg_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_request/$exit
      -- CP-element group 48: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_request/ack
      -- 
    ack_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_351_final_reg_ack_0, ack => zeropad3D_CP_676_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	583 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	82 
    -- CP-element group 49:  members (19) 
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_base_plus_offset/sum_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_base_addr_resize/base_resize_req
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_base_plus_offset/sum_rename_req
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_word_addrgen/$entry
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_word_addrgen/$exit
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_word_addrgen/root_register_req
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_word_addrgen/root_register_ack
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_base_plus_offset/$exit
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_base_addr_resize/base_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_base_plus_offset/$entry
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_base_addr_resize/$exit
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_base_addr_resize/$entry
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_base_address_resized
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_root_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_word_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_base_address_calculated
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_complete/$exit
      -- CP-element group 49: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_complete/ack
      -- 
    ack_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_351_final_reg_ack_1, ack => zeropad3D_CP_676_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	583 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_update_start_
      -- CP-element group 50: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_Update/cr
      -- 
    ra_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_354_inst_ack_0, ack => zeropad3D_CP_676_elements(50)); -- 
    cr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(50), ack => RPIPE_zeropad_input_pipe_354_inst_req_1); -- 
    -- CP-element group 51:  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	54 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_Sample/rr
      -- 
    ca_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_354_inst_ack_1, ack => zeropad3D_CP_676_elements(51)); -- 
    rr_1380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(51), ack => type_cast_358_inst_req_0); -- 
    rr_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(51), ack => RPIPE_zeropad_input_pipe_367_inst_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_Sample/ra
      -- 
    ra_1381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_0, ack => zeropad3D_CP_676_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	583 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	82 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_Update/ca
      -- 
    ca_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_1, ack => zeropad3D_CP_676_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_update_start_
      -- CP-element group 54: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_Update/cr
      -- 
    ra_1395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_367_inst_ack_0, ack => zeropad3D_CP_676_elements(54)); -- 
    cr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(54), ack => RPIPE_zeropad_input_pipe_367_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_367_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_Sample/rr
      -- 
    ca_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_367_inst_ack_1, ack => zeropad3D_CP_676_elements(55)); -- 
    rr_1408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(55), ack => type_cast_371_inst_req_0); -- 
    rr_1422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(55), ack => RPIPE_zeropad_input_pipe_385_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_Sample/ra
      -- 
    ra_1409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_0, ack => zeropad3D_CP_676_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	583 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	82 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_Update/ca
      -- 
    ca_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_1, ack => zeropad3D_CP_676_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_update_start_
      -- CP-element group 58: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_Update/cr
      -- 
    ra_1423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_385_inst_ack_0, ack => zeropad3D_CP_676_elements(58)); -- 
    cr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(58), ack => RPIPE_zeropad_input_pipe_385_inst_req_1); -- 
    -- CP-element group 59:  fork  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	62 
    -- CP-element group 59:  members (9) 
      -- CP-element group 59: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_385_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_Sample/rr
      -- 
    ca_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_385_inst_ack_1, ack => zeropad3D_CP_676_elements(59)); -- 
    rr_1436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(59), ack => type_cast_389_inst_req_0); -- 
    rr_1450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(59), ack => RPIPE_zeropad_input_pipe_403_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_Sample/ra
      -- 
    ra_1437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_389_inst_ack_0, ack => zeropad3D_CP_676_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	583 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	82 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_Update/ca
      -- 
    ca_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_389_inst_ack_1, ack => zeropad3D_CP_676_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_update_start_
      -- CP-element group 62: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_Update/cr
      -- 
    ra_1451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_403_inst_ack_0, ack => zeropad3D_CP_676_elements(62)); -- 
    cr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(62), ack => RPIPE_zeropad_input_pipe_403_inst_req_1); -- 
    -- CP-element group 63:  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_403_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_Sample/rr
      -- 
    ca_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_403_inst_ack_1, ack => zeropad3D_CP_676_elements(63)); -- 
    rr_1464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(63), ack => type_cast_407_inst_req_0); -- 
    rr_1478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(63), ack => RPIPE_zeropad_input_pipe_421_inst_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_Sample/ra
      -- 
    ra_1465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_407_inst_ack_0, ack => zeropad3D_CP_676_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	583 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	82 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_Update/ca
      -- 
    ca_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_407_inst_ack_1, ack => zeropad3D_CP_676_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_update_start_
      -- CP-element group 66: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_Update/cr
      -- 
    ra_1479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_421_inst_ack_0, ack => zeropad3D_CP_676_elements(66)); -- 
    cr_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(66), ack => RPIPE_zeropad_input_pipe_421_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	70 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_421_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_Sample/rr
      -- 
    ca_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_421_inst_ack_1, ack => zeropad3D_CP_676_elements(67)); -- 
    rr_1492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(67), ack => type_cast_425_inst_req_0); -- 
    rr_1506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(67), ack => RPIPE_zeropad_input_pipe_439_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_Sample/ra
      -- 
    ra_1493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_425_inst_ack_0, ack => zeropad3D_CP_676_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	583 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	82 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_Update/ca
      -- CP-element group 69: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_update_completed_
      -- 
    ca_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_425_inst_ack_1, ack => zeropad3D_CP_676_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_update_start_
      -- CP-element group 70: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_Update/cr
      -- 
    ra_1507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_439_inst_ack_0, ack => zeropad3D_CP_676_elements(70)); -- 
    cr_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(70), ack => RPIPE_zeropad_input_pipe_439_inst_req_1); -- 
    -- CP-element group 71:  fork  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: 	74 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_439_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_Sample/$entry
      -- 
    ca_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_439_inst_ack_1, ack => zeropad3D_CP_676_elements(71)); -- 
    rr_1534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(71), ack => RPIPE_zeropad_input_pipe_457_inst_req_0); -- 
    rr_1520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(71), ack => type_cast_443_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_Sample/$exit
      -- 
    ra_1521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_0, ack => zeropad3D_CP_676_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	583 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	82 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_update_completed_
      -- 
    ca_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_1, ack => zeropad3D_CP_676_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	71 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_update_start_
      -- CP-element group 74: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_sample_completed_
      -- 
    ra_1535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_457_inst_ack_0, ack => zeropad3D_CP_676_elements(74)); -- 
    cr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(74), ack => RPIPE_zeropad_input_pipe_457_inst_req_1); -- 
    -- CP-element group 75:  fork  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (9) 
      -- CP-element group 75: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_457_update_completed_
      -- 
    ca_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_457_inst_ack_1, ack => zeropad3D_CP_676_elements(75)); -- 
    rr_1548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(75), ack => type_cast_461_inst_req_0); -- 
    rr_1562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(75), ack => RPIPE_zeropad_input_pipe_475_inst_req_0); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_sample_completed_
      -- 
    ra_1549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_0, ack => zeropad3D_CP_676_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	583 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	82 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_Update/$exit
      -- 
    ca_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_1, ack => zeropad3D_CP_676_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_update_start_
      -- CP-element group 78: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_Update/cr
      -- 
    ra_1563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_475_inst_ack_0, ack => zeropad3D_CP_676_elements(78)); -- 
    cr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(78), ack => RPIPE_zeropad_input_pipe_475_inst_req_1); -- 
    -- CP-element group 79:  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (6) 
      -- CP-element group 79: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_475_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_Sample/rr
      -- 
    ca_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_475_inst_ack_1, ack => zeropad3D_CP_676_elements(79)); -- 
    rr_1576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(79), ack => type_cast_479_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_Sample/ra
      -- 
    ra_1577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_479_inst_ack_0, ack => zeropad3D_CP_676_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	583 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_Update/$exit
      -- 
    ca_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_479_inst_ack_1, ack => zeropad3D_CP_676_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	73 
    -- CP-element group 82: 	49 
    -- CP-element group 82: 	53 
    -- CP-element group 82: 	57 
    -- CP-element group 82: 	61 
    -- CP-element group 82: 	65 
    -- CP-element group 82: 	69 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (9) 
      -- CP-element group 82: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/ptr_deref_487_Split/split_req
      -- CP-element group 82: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/ptr_deref_487_Split/$entry
      -- CP-element group 82: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/ptr_deref_487_Split/$exit
      -- CP-element group 82: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/ptr_deref_487_Split/split_ack
      -- CP-element group 82: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/word_access_start/$entry
      -- CP-element group 82: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/word_access_start/word_0/$entry
      -- CP-element group 82: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/word_access_start/word_0/rr
      -- CP-element group 82: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_sample_start_
      -- 
    rr_1620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(82), ack => ptr_deref_487_store_0_req_0); -- 
    zeropad3D_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(73) & zeropad3D_CP_676_elements(49) & zeropad3D_CP_676_elements(53) & zeropad3D_CP_676_elements(57) & zeropad3D_CP_676_elements(61) & zeropad3D_CP_676_elements(65) & zeropad3D_CP_676_elements(69) & zeropad3D_CP_676_elements(77) & zeropad3D_CP_676_elements(81);
      gj_zeropad3D_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/word_access_start/$exit
      -- CP-element group 83: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/word_access_start/word_0/ra
      -- CP-element group 83: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Sample/word_access_start/word_0/$exit
      -- 
    ra_1621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_487_store_0_ack_0, ack => zeropad3D_CP_676_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	583 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Update/word_access_complete/word_0/ca
      -- CP-element group 84: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Update/word_access_complete/word_0/$exit
      -- CP-element group 84: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Update/word_access_complete/$exit
      -- CP-element group 84: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_update_completed_
      -- 
    ca_1632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_487_store_0_ack_1, ack => zeropad3D_CP_676_elements(84)); -- 
    -- CP-element group 85:  branch  join  transition  place  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	46 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (10) 
      -- CP-element group 85: 	 branch_block_stmt_223/if_stmt_501_else_link/$entry
      -- CP-element group 85: 	 branch_block_stmt_223/if_stmt_501_eval_test/$exit
      -- CP-element group 85: 	 branch_block_stmt_223/if_stmt_501__entry__
      -- CP-element group 85: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500__exit__
      -- CP-element group 85: 	 branch_block_stmt_223/if_stmt_501_eval_test/$entry
      -- CP-element group 85: 	 branch_block_stmt_223/if_stmt_501_dead_link/$entry
      -- CP-element group 85: 	 branch_block_stmt_223/if_stmt_501_eval_test/branch_req
      -- CP-element group 85: 	 branch_block_stmt_223/if_stmt_501_if_link/$entry
      -- CP-element group 85: 	 branch_block_stmt_223/R_exitcond8_502_place
      -- CP-element group 85: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/$exit
      -- 
    branch_req_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(85), ack => if_stmt_501_branch_req_0); -- 
    zeropad3D_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(46) & zeropad3D_CP_676_elements(84);
      gj_zeropad3D_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  merge  transition  place  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	584 
    -- CP-element group 86:  members (13) 
      -- CP-element group 86: 	 branch_block_stmt_223/merge_stmt_507__exit__
      -- CP-element group 86: 	 branch_block_stmt_223/forx_xendx_xloopexit_forx_xend
      -- CP-element group 86: 	 branch_block_stmt_223/if_stmt_501_if_link/$exit
      -- CP-element group 86: 	 branch_block_stmt_223/if_stmt_501_if_link/if_choice_transition
      -- CP-element group 86: 	 branch_block_stmt_223/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 86: 	 branch_block_stmt_223/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_223/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_223/merge_stmt_507_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_223/merge_stmt_507_PhiAck/$entry
      -- CP-element group 86: 	 branch_block_stmt_223/merge_stmt_507_PhiAck/$exit
      -- CP-element group 86: 	 branch_block_stmt_223/merge_stmt_507_PhiAck/dummy
      -- CP-element group 86: 	 branch_block_stmt_223/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_223/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_501_branch_ack_1, ack => zeropad3D_CP_676_elements(86)); -- 
    -- CP-element group 87:  fork  transition  place  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	579 
    -- CP-element group 87: 	580 
    -- CP-element group 87:  members (12) 
      -- CP-element group 87: 	 branch_block_stmt_223/if_stmt_501_else_link/$exit
      -- CP-element group 87: 	 branch_block_stmt_223/if_stmt_501_else_link/else_choice_transition
      -- CP-element group 87: 	 branch_block_stmt_223/forx_xbody_forx_xbody
      -- CP-element group 87: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 87: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/$entry
      -- CP-element group 87: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/$entry
      -- CP-element group 87: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/$entry
      -- CP-element group 87: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/SplitProtocol/$entry
      -- CP-element group 87: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/SplitProtocol/Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/SplitProtocol/Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/SplitProtocol/Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_501_branch_ack_0, ack => zeropad3D_CP_676_elements(87)); -- 
    rr_6674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(87), ack => type_cast_344_inst_req_0); -- 
    cr_6679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(87), ack => type_cast_344_inst_req_1); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	584 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Sample/word_access_start/$exit
      -- CP-element group 88: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Sample/word_access_start/word_0/$exit
      -- CP-element group 88: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Sample/word_access_start/word_0/ra
      -- CP-element group 88: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Sample/$exit
      -- 
    ra_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_512_load_0_ack_0, ack => zeropad3D_CP_676_elements(88)); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	584 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	98 
    -- CP-element group 89:  members (12) 
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/word_access_complete/$exit
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/LOAD_pad_512_Merge/merge_ack
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/LOAD_pad_512_Merge/merge_req
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/LOAD_pad_512_Merge/$exit
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/LOAD_pad_512_Merge/$entry
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/word_access_complete/word_0/ca
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/word_access_complete/word_0/$exit
      -- 
    ca_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_512_load_0_ack_1, ack => zeropad3D_CP_676_elements(89)); -- 
    rr_1751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(89), ack => type_cast_537_inst_req_0); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	584 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_sample_completed_
      -- 
    ra_1696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_516_inst_ack_0, ack => zeropad3D_CP_676_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	584 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	104 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_update_completed_
      -- 
    ca_1701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_516_inst_ack_1, ack => zeropad3D_CP_676_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	584 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_sample_completed_
      -- 
    ra_1710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_0, ack => zeropad3D_CP_676_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	584 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	104 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_Update/ca
      -- CP-element group 93: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_update_completed_
      -- 
    ca_1715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_1, ack => zeropad3D_CP_676_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	584 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_Sample/ra
      -- 
    ra_1724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_524_inst_ack_0, ack => zeropad3D_CP_676_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	584 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	104 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_Update/$exit
      -- 
    ca_1729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_524_inst_ack_1, ack => zeropad3D_CP_676_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	584 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_sample_completed_
      -- 
    ra_1738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_528_inst_ack_0, ack => zeropad3D_CP_676_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	584 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	104 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_Update/ca
      -- 
    ca_1743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_528_inst_ack_1, ack => zeropad3D_CP_676_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	89 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_Sample/$exit
      -- 
    ra_1752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_537_inst_ack_0, ack => zeropad3D_CP_676_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	584 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	104 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_update_completed_
      -- 
    ca_1757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_537_inst_ack_1, ack => zeropad3D_CP_676_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	584 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_sample_completed_
      -- 
    ra_1766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_0, ack => zeropad3D_CP_676_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	584 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_update_completed_
      -- 
    ca_1771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_541_inst_ack_1, ack => zeropad3D_CP_676_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	584 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_sample_completed_
      -- 
    ra_1780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_0, ack => zeropad3D_CP_676_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	584 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_update_completed_
      -- 
    ca_1785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_1, ack => zeropad3D_CP_676_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	91 
    -- CP-element group 104: 	93 
    -- CP-element group 104: 	95 
    -- CP-element group 104: 	97 
    -- CP-element group 104: 	99 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	585 
    -- CP-element group 104: 	586 
    -- CP-element group 104: 	587 
    -- CP-element group 104:  members (10) 
      -- CP-element group 104: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/$exit
      -- CP-element group 104: 	 branch_block_stmt_223/forx_xend_whilex_xbody
      -- CP-element group 104: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619__exit__
      -- CP-element group 104: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/$entry
      -- CP-element group 104: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_622/$entry
      -- CP-element group 104: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_630/$entry
      -- CP-element group 104: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_637/$entry
      -- CP-element group 104: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/$entry
      -- 
    zeropad3D_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(91) & zeropad3D_CP_676_elements(93) & zeropad3D_CP_676_elements(95) & zeropad3D_CP_676_elements(97) & zeropad3D_CP_676_elements(99) & zeropad3D_CP_676_elements(101) & zeropad3D_CP_676_elements(103);
      gj_zeropad3D_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	603 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_sample_completed_
      -- 
    ra_1797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_648_inst_ack_0, ack => zeropad3D_CP_676_elements(105)); -- 
    -- CP-element group 106:  branch  transition  place  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	603 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (13) 
      -- CP-element group 106: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674__exit__
      -- CP-element group 106: 	 branch_block_stmt_223/if_stmt_675_eval_test/$entry
      -- CP-element group 106: 	 branch_block_stmt_223/if_stmt_675_eval_test/$exit
      -- CP-element group 106: 	 branch_block_stmt_223/if_stmt_675__entry__
      -- CP-element group 106: 	 branch_block_stmt_223/if_stmt_675_eval_test/branch_req
      -- CP-element group 106: 	 branch_block_stmt_223/if_stmt_675_dead_link/$entry
      -- CP-element group 106: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/$exit
      -- CP-element group 106: 	 branch_block_stmt_223/if_stmt_675_else_link/$entry
      -- CP-element group 106: 	 branch_block_stmt_223/if_stmt_675_if_link/$entry
      -- CP-element group 106: 	 branch_block_stmt_223/R_orx_xcond_676_place
      -- 
    ca_1802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_648_inst_ack_1, ack => zeropad3D_CP_676_elements(106)); -- 
    branch_req_1810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(106), ack => if_stmt_675_branch_req_0); -- 
    -- CP-element group 107:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (18) 
      -- CP-element group 107: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_Update/cr
      -- CP-element group 107: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711__entry__
      -- CP-element group 107: 	 branch_block_stmt_223/merge_stmt_681__exit__
      -- CP-element group 107: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_update_start_
      -- CP-element group 107: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/$entry
      -- CP-element group 107: 	 branch_block_stmt_223/whilex_xbody_lorx_xlhsx_xfalse122
      -- CP-element group 107: 	 branch_block_stmt_223/if_stmt_675_if_link/if_choice_transition
      -- CP-element group 107: 	 branch_block_stmt_223/if_stmt_675_if_link/$exit
      -- CP-element group 107: 	 branch_block_stmt_223/whilex_xbody_lorx_xlhsx_xfalse122_PhiReq/$entry
      -- CP-element group 107: 	 branch_block_stmt_223/whilex_xbody_lorx_xlhsx_xfalse122_PhiReq/$exit
      -- CP-element group 107: 	 branch_block_stmt_223/merge_stmt_681_PhiReqMerge
      -- CP-element group 107: 	 branch_block_stmt_223/merge_stmt_681_PhiAck/$entry
      -- CP-element group 107: 	 branch_block_stmt_223/merge_stmt_681_PhiAck/$exit
      -- CP-element group 107: 	 branch_block_stmt_223/merge_stmt_681_PhiAck/dummy
      -- 
    if_choice_transition_1815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_675_branch_ack_1, ack => zeropad3D_CP_676_elements(107)); -- 
    cr_1837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(107), ack => type_cast_685_inst_req_1); -- 
    rr_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(107), ack => type_cast_685_inst_req_0); -- 
    -- CP-element group 108:  transition  place  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	604 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_223/whilex_xbody_ifx_xthen
      -- CP-element group 108: 	 branch_block_stmt_223/if_stmt_675_else_link/else_choice_transition
      -- CP-element group 108: 	 branch_block_stmt_223/if_stmt_675_else_link/$exit
      -- CP-element group 108: 	 branch_block_stmt_223/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 108: 	 branch_block_stmt_223/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_1819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_675_branch_ack_0, ack => zeropad3D_CP_676_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_sample_completed_
      -- 
    ra_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_685_inst_ack_0, ack => zeropad3D_CP_676_elements(109)); -- 
    -- CP-element group 110:  branch  transition  place  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (13) 
      -- CP-element group 110: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_223/if_stmt_712__entry__
      -- CP-element group 110: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711__exit__
      -- CP-element group 110: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_Update/ca
      -- CP-element group 110: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/type_cast_685_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_223/if_stmt_712_else_link/$entry
      -- CP-element group 110: 	 branch_block_stmt_223/if_stmt_712_if_link/$entry
      -- CP-element group 110: 	 branch_block_stmt_223/R_orx_xcond1849_713_place
      -- CP-element group 110: 	 branch_block_stmt_223/if_stmt_712_eval_test/branch_req
      -- CP-element group 110: 	 branch_block_stmt_223/if_stmt_712_eval_test/$exit
      -- CP-element group 110: 	 branch_block_stmt_223/if_stmt_712_eval_test/$entry
      -- CP-element group 110: 	 branch_block_stmt_223/assign_stmt_686_to_assign_stmt_711/$exit
      -- CP-element group 110: 	 branch_block_stmt_223/if_stmt_712_dead_link/$entry
      -- 
    ca_1838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_685_inst_ack_1, ack => zeropad3D_CP_676_elements(110)); -- 
    branch_req_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(110), ack => if_stmt_712_branch_req_0); -- 
    -- CP-element group 111:  fork  transition  place  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	127 
    -- CP-element group 111: 	128 
    -- CP-element group 111: 	130 
    -- CP-element group 111: 	132 
    -- CP-element group 111: 	134 
    -- CP-element group 111: 	136 
    -- CP-element group 111: 	138 
    -- CP-element group 111: 	140 
    -- CP-element group 111: 	142 
    -- CP-element group 111: 	145 
    -- CP-element group 111:  members (46) 
      -- CP-element group 111: 	 branch_block_stmt_223/lorx_xlhsx_xfalse122_ifx_xelse
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882__entry__
      -- CP-element group 111: 	 branch_block_stmt_223/merge_stmt_777__exit__
      -- CP-element group 111: 	 branch_block_stmt_223/if_stmt_712_if_link/if_choice_transition
      -- CP-element group 111: 	 branch_block_stmt_223/if_stmt_712_if_link/$exit
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_update_start_
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_update_start_
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_update_start_
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_final_index_sum_regn_update_start
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_final_index_sum_regn_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_final_index_sum_regn_Update/req
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_complete/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_complete/req
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_update_start_
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/word_access_complete/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/word_access_complete/word_0/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/word_access_complete/word_0/cr
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_update_start_
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_update_start_
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_final_index_sum_regn_update_start
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_final_index_sum_regn_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_final_index_sum_regn_Update/req
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_complete/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_complete/req
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_update_start_
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Update/word_access_complete/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Update/word_access_complete/word_0/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Update/word_access_complete/word_0/cr
      -- CP-element group 111: 	 branch_block_stmt_223/lorx_xlhsx_xfalse122_ifx_xelse_PhiReq/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/lorx_xlhsx_xfalse122_ifx_xelse_PhiReq/$exit
      -- CP-element group 111: 	 branch_block_stmt_223/merge_stmt_777_PhiReqMerge
      -- CP-element group 111: 	 branch_block_stmt_223/merge_stmt_777_PhiAck/$entry
      -- CP-element group 111: 	 branch_block_stmt_223/merge_stmt_777_PhiAck/$exit
      -- CP-element group 111: 	 branch_block_stmt_223/merge_stmt_777_PhiAck/dummy
      -- 
    if_choice_transition_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_712_branch_ack_1, ack => zeropad3D_CP_676_elements(111)); -- 
    rr_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => type_cast_781_inst_req_0); -- 
    cr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => type_cast_781_inst_req_1); -- 
    cr_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => type_cast_845_inst_req_1); -- 
    req_2059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => array_obj_ref_851_index_offset_req_1); -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => addr_of_852_final_reg_req_1); -- 
    cr_2119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => ptr_deref_856_load_0_req_1); -- 
    cr_2138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => type_cast_870_inst_req_1); -- 
    req_2169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => array_obj_ref_876_index_offset_req_1); -- 
    req_2184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => addr_of_877_final_reg_req_1); -- 
    cr_2234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => ptr_deref_880_store_0_req_1); -- 
    -- CP-element group 112:  transition  place  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	604 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_223/lorx_xlhsx_xfalse122_ifx_xthen
      -- CP-element group 112: 	 branch_block_stmt_223/if_stmt_712_else_link/else_choice_transition
      -- CP-element group 112: 	 branch_block_stmt_223/if_stmt_712_else_link/$exit
      -- CP-element group 112: 	 branch_block_stmt_223/lorx_xlhsx_xfalse122_ifx_xthen_PhiReq/$entry
      -- CP-element group 112: 	 branch_block_stmt_223/lorx_xlhsx_xfalse122_ifx_xthen_PhiReq/$exit
      -- 
    else_choice_transition_1855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_712_branch_ack_0, ack => zeropad3D_CP_676_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	604 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_Sample/$exit
      -- 
    ra_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_0, ack => zeropad3D_CP_676_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	604 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	117 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_Update/ca
      -- 
    ca_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_722_inst_ack_1, ack => zeropad3D_CP_676_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	604 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_sample_completed_
      -- 
    ra_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_0, ack => zeropad3D_CP_676_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	604 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_update_completed_
      -- 
    ca_1888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_727_inst_ack_1, ack => zeropad3D_CP_676_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	114 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_Sample/$entry
      -- 
    rr_1896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(117), ack => type_cast_762_inst_req_0); -- 
    zeropad3D_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(114) & zeropad3D_CP_676_elements(116);
      gj_zeropad3D_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_Sample/ra
      -- CP-element group 118: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_Sample/$exit
      -- 
    ra_1897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_762_inst_ack_0, ack => zeropad3D_CP_676_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	604 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (16) 
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_scale_1/$entry
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_scale_1/$exit
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_scale_1/scale_rename_req
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_scale_1/scale_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_final_index_sum_regn_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_resize_1/index_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_resize_1/index_resize_req
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_resize_1/$exit
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_resize_1/$entry
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_computed_1
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_scaled_1
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_index_resized_1
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_final_index_sum_regn_Sample/req
      -- CP-element group 119: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_Update/ca
      -- 
    ca_1902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_762_inst_ack_1, ack => zeropad3D_CP_676_elements(119)); -- 
    req_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(119), ack => array_obj_ref_768_index_offset_req_0); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	126 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_final_index_sum_regn_sample_complete
      -- CP-element group 120: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_final_index_sum_regn_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_final_index_sum_regn_Sample/ack
      -- 
    ack_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_768_index_offset_ack_0, ack => zeropad3D_CP_676_elements(120)); -- 
    -- CP-element group 121:  transition  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	604 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (11) 
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_request/$entry
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_request/req
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_base_plus_offset/sum_rename_ack
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_offset_calculated
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_root_address_calculated
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_base_plus_offset/sum_rename_req
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_base_plus_offset/$exit
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_base_plus_offset/$entry
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_final_index_sum_regn_Update/ack
      -- CP-element group 121: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_final_index_sum_regn_Update/$exit
      -- 
    ack_1933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_768_index_offset_ack_1, ack => zeropad3D_CP_676_elements(121)); -- 
    req_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(121), ack => addr_of_769_final_reg_req_0); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_request/$exit
      -- CP-element group 122: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_request/ack
      -- CP-element group 122: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_sample_completed_
      -- 
    ack_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_769_final_reg_ack_0, ack => zeropad3D_CP_676_elements(122)); -- 
    -- CP-element group 123:  join  fork  transition  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	604 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (28) 
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_word_addrgen/$exit
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_word_addrgen/$entry
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_base_addr_resize/base_resize_ack
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_complete/ack
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/ptr_deref_772_Split/split_ack
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_complete/$exit
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/ptr_deref_772_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_base_addr_resize/base_resize_req
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_base_addr_resize/$exit
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/ptr_deref_772_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/ptr_deref_772_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_base_addr_resize/$entry
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_base_address_resized
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_base_plus_offset/sum_rename_ack
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_base_plus_offset/sum_rename_req
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_root_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_word_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_base_plus_offset/$exit
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_word_addrgen/root_register_ack
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_base_plus_offset/$entry
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/word_access_start/word_0/rr
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_base_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_word_addrgen/root_register_req
      -- 
    ack_1948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_769_final_reg_ack_1, ack => zeropad3D_CP_676_elements(123)); -- 
    rr_1986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(123), ack => ptr_deref_772_store_0_req_0); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/word_access_start/word_0/ra
      -- CP-element group 124: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Sample/word_access_start/word_0/$exit
      -- 
    ra_1987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_772_store_0_ack_0, ack => zeropad3D_CP_676_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	604 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Update/word_access_complete/word_0/ca
      -- 
    ca_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_772_store_0_ack_1, ack => zeropad3D_CP_676_elements(125)); -- 
    -- CP-element group 126:  join  transition  place  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	120 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	605 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775__exit__
      -- CP-element group 126: 	 branch_block_stmt_223/ifx_xthen_ifx_xend
      -- CP-element group 126: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/$exit
      -- CP-element group 126: 	 branch_block_stmt_223/ifx_xthen_ifx_xend_PhiReq/$entry
      -- CP-element group 126: 	 branch_block_stmt_223/ifx_xthen_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(120) & zeropad3D_CP_676_elements(125);
      gj_zeropad3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	111 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_Sample/ra
      -- 
    ra_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_0, ack => zeropad3D_CP_676_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	111 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128: 	137 
    -- CP-element group 128:  members (9) 
      -- CP-element group 128: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_781_Update/ca
      -- CP-element group 128: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_Sample/rr
      -- 
    ca_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_781_inst_ack_1, ack => zeropad3D_CP_676_elements(128)); -- 
    rr_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => type_cast_845_inst_req_0); -- 
    rr_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => type_cast_870_inst_req_0); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_Sample/ra
      -- 
    ra_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_845_inst_ack_0, ack => zeropad3D_CP_676_elements(129)); -- 
    -- CP-element group 130:  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	111 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (16) 
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_845_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_resized_1
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_scaled_1
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_computed_1
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_resize_1/$entry
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_resize_1/$exit
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_resize_1/index_resize_req
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_resize_1/index_resize_ack
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_scale_1/$entry
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_scale_1/$exit
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_scale_1/scale_rename_req
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_index_scale_1/scale_rename_ack
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_final_index_sum_regn_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_final_index_sum_regn_Sample/req
      -- 
    ca_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_845_inst_ack_1, ack => zeropad3D_CP_676_elements(130)); -- 
    req_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(130), ack => array_obj_ref_851_index_offset_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	146 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_final_index_sum_regn_sample_complete
      -- CP-element group 131: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_final_index_sum_regn_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_final_index_sum_regn_Sample/ack
      -- 
    ack_2055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_851_index_offset_ack_0, ack => zeropad3D_CP_676_elements(131)); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	111 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (11) 
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_root_address_calculated
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_offset_calculated
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_final_index_sum_regn_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_final_index_sum_regn_Update/ack
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_base_plus_offset/$entry
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_base_plus_offset/$exit
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_base_plus_offset/sum_rename_req
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_851_base_plus_offset/sum_rename_ack
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_request/$entry
      -- CP-element group 132: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_request/req
      -- 
    ack_2060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_851_index_offset_ack_1, ack => zeropad3D_CP_676_elements(132)); -- 
    req_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(132), ack => addr_of_852_final_reg_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_request/$exit
      -- CP-element group 133: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_request/ack
      -- 
    ack_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_852_final_reg_ack_0, ack => zeropad3D_CP_676_elements(133)); -- 
    -- CP-element group 134:  join  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	111 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (24) 
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_complete/$exit
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_852_complete/ack
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_base_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_word_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_root_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_base_address_resized
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_base_addr_resize/$entry
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_base_addr_resize/$exit
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_base_addr_resize/base_resize_req
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_base_addr_resize/base_resize_ack
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_base_plus_offset/$entry
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_base_plus_offset/$exit
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_base_plus_offset/sum_rename_req
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_base_plus_offset/sum_rename_ack
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_word_addrgen/$entry
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_word_addrgen/$exit
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_word_addrgen/root_register_req
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_word_addrgen/root_register_ack
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Sample/word_access_start/$entry
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Sample/word_access_start/word_0/$entry
      -- CP-element group 134: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Sample/word_access_start/word_0/rr
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_852_final_reg_ack_1, ack => zeropad3D_CP_676_elements(134)); -- 
    rr_2108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(134), ack => ptr_deref_856_load_0_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (5) 
      -- CP-element group 135: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Sample/word_access_start/$exit
      -- CP-element group 135: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Sample/word_access_start/word_0/$exit
      -- CP-element group 135: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Sample/word_access_start/word_0/ra
      -- 
    ra_2109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_856_load_0_ack_0, ack => zeropad3D_CP_676_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	111 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	143 
    -- CP-element group 136:  members (9) 
      -- CP-element group 136: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/word_access_complete/$exit
      -- CP-element group 136: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/word_access_complete/word_0/$exit
      -- CP-element group 136: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/word_access_complete/word_0/ca
      -- CP-element group 136: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/ptr_deref_856_Merge/$entry
      -- CP-element group 136: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/ptr_deref_856_Merge/$exit
      -- CP-element group 136: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/ptr_deref_856_Merge/merge_req
      -- CP-element group 136: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_856_Update/ptr_deref_856_Merge/merge_ack
      -- 
    ca_2120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_856_load_0_ack_1, ack => zeropad3D_CP_676_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	128 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_Sample/ra
      -- 
    ra_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_870_inst_ack_0, ack => zeropad3D_CP_676_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	111 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (16) 
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/type_cast_870_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_resized_1
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_scaled_1
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_computed_1
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_resize_1/$entry
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_resize_1/$exit
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_resize_1/index_resize_req
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_resize_1/index_resize_ack
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_scale_1/$entry
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_scale_1/$exit
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_scale_1/scale_rename_req
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_index_scale_1/scale_rename_ack
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_final_index_sum_regn_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_final_index_sum_regn_Sample/req
      -- 
    ca_2139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_870_inst_ack_1, ack => zeropad3D_CP_676_elements(138)); -- 
    req_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(138), ack => array_obj_ref_876_index_offset_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	146 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_final_index_sum_regn_sample_complete
      -- CP-element group 139: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_final_index_sum_regn_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_final_index_sum_regn_Sample/ack
      -- 
    ack_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_876_index_offset_ack_0, ack => zeropad3D_CP_676_elements(139)); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	111 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (11) 
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_root_address_calculated
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_offset_calculated
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_final_index_sum_regn_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_final_index_sum_regn_Update/ack
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_base_plus_offset/$entry
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_base_plus_offset/$exit
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_base_plus_offset/sum_rename_req
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/array_obj_ref_876_base_plus_offset/sum_rename_ack
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_request/$entry
      -- CP-element group 140: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_request/req
      -- 
    ack_2170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_876_index_offset_ack_1, ack => zeropad3D_CP_676_elements(140)); -- 
    req_2179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(140), ack => addr_of_877_final_reg_req_0); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_request/$exit
      -- CP-element group 141: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_request/ack
      -- 
    ack_2180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_877_final_reg_ack_0, ack => zeropad3D_CP_676_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	111 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (19) 
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_complete/$exit
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/addr_of_877_complete/ack
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_base_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_word_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_root_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_base_address_resized
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_base_addr_resize/$entry
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_base_addr_resize/$exit
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_base_addr_resize/base_resize_req
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_base_addr_resize/base_resize_ack
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_base_plus_offset/$entry
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_base_plus_offset/$exit
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_base_plus_offset/sum_rename_req
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_base_plus_offset/sum_rename_ack
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_word_addrgen/$entry
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_word_addrgen/$exit
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_word_addrgen/root_register_req
      -- CP-element group 142: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_word_addrgen/root_register_ack
      -- 
    ack_2185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_877_final_reg_ack_1, ack => zeropad3D_CP_676_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	136 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (9) 
      -- CP-element group 143: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/ptr_deref_880_Split/$entry
      -- CP-element group 143: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/ptr_deref_880_Split/$exit
      -- CP-element group 143: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/ptr_deref_880_Split/split_req
      -- CP-element group 143: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/ptr_deref_880_Split/split_ack
      -- CP-element group 143: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/word_access_start/word_0/rr
      -- 
    rr_2223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(143), ack => ptr_deref_880_store_0_req_0); -- 
    zeropad3D_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(136) & zeropad3D_CP_676_elements(142);
      gj_zeropad3D_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Sample/word_access_start/word_0/ra
      -- 
    ra_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_880_store_0_ack_0, ack => zeropad3D_CP_676_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	111 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/ptr_deref_880_Update/word_access_complete/word_0/ca
      -- 
    ca_2235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_880_store_0_ack_1, ack => zeropad3D_CP_676_elements(145)); -- 
    -- CP-element group 146:  join  transition  place  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	131 
    -- CP-element group 146: 	139 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	605 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882__exit__
      -- CP-element group 146: 	 branch_block_stmt_223/ifx_xelse_ifx_xend
      -- CP-element group 146: 	 branch_block_stmt_223/assign_stmt_782_to_assign_stmt_882/$exit
      -- CP-element group 146: 	 branch_block_stmt_223/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 146: 	 branch_block_stmt_223/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(131) & zeropad3D_CP_676_elements(139) & zeropad3D_CP_676_elements(145);
      gj_zeropad3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	605 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_Sample/ra
      -- 
    ra_2247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_888_inst_ack_0, ack => zeropad3D_CP_676_elements(147)); -- 
    -- CP-element group 148:  branch  transition  place  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	605 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (13) 
      -- CP-element group 148: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902__exit__
      -- CP-element group 148: 	 branch_block_stmt_223/if_stmt_903__entry__
      -- CP-element group 148: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/$exit
      -- CP-element group 148: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_223/if_stmt_903_dead_link/$entry
      -- CP-element group 148: 	 branch_block_stmt_223/if_stmt_903_eval_test/$entry
      -- CP-element group 148: 	 branch_block_stmt_223/if_stmt_903_eval_test/$exit
      -- CP-element group 148: 	 branch_block_stmt_223/if_stmt_903_eval_test/branch_req
      -- CP-element group 148: 	 branch_block_stmt_223/R_cmp210_904_place
      -- CP-element group 148: 	 branch_block_stmt_223/if_stmt_903_if_link/$entry
      -- CP-element group 148: 	 branch_block_stmt_223/if_stmt_903_else_link/$entry
      -- 
    ca_2252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_888_inst_ack_1, ack => zeropad3D_CP_676_elements(148)); -- 
    branch_req_2260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(148), ack => if_stmt_903_branch_req_0); -- 
    -- CP-element group 149:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	614 
    -- CP-element group 149: 	615 
    -- CP-element group 149: 	617 
    -- CP-element group 149: 	618 
    -- CP-element group 149: 	620 
    -- CP-element group 149: 	621 
    -- CP-element group 149:  members (40) 
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253
      -- CP-element group 149: 	 branch_block_stmt_223/assign_stmt_915__exit__
      -- CP-element group 149: 	 branch_block_stmt_223/assign_stmt_915__entry__
      -- CP-element group 149: 	 branch_block_stmt_223/merge_stmt_909__exit__
      -- CP-element group 149: 	 branch_block_stmt_223/if_stmt_903_if_link/$exit
      -- CP-element group 149: 	 branch_block_stmt_223/if_stmt_903_if_link/if_choice_transition
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xend_ifx_xthen212
      -- CP-element group 149: 	 branch_block_stmt_223/assign_stmt_915/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/assign_stmt_915/$exit
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/SplitProtocol/Update/cr
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/SplitProtocol/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/SplitProtocol/Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/SplitProtocol/Sample/rr
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/SplitProtocol/Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/SplitProtocol/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/SplitProtocol/Update/cr
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/SplitProtocol/Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/SplitProtocol/Sample/rr
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/SplitProtocol/Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/SplitProtocol/Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/SplitProtocol/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/SplitProtocol/Sample/rr
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/SplitProtocol/Update/cr
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/SplitProtocol/Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xend_ifx_xthen212_PhiReq/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/ifx_xend_ifx_xthen212_PhiReq/$exit
      -- CP-element group 149: 	 branch_block_stmt_223/merge_stmt_909_PhiReqMerge
      -- CP-element group 149: 	 branch_block_stmt_223/merge_stmt_909_PhiAck/$entry
      -- CP-element group 149: 	 branch_block_stmt_223/merge_stmt_909_PhiAck/$exit
      -- CP-element group 149: 	 branch_block_stmt_223/merge_stmt_909_PhiAck/dummy
      -- 
    if_choice_transition_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_903_branch_ack_1, ack => zeropad3D_CP_676_elements(149)); -- 
    cr_6989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(149), ack => type_cast_976_inst_req_1); -- 
    rr_6961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(149), ack => type_cast_970_inst_req_0); -- 
    cr_7012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(149), ack => type_cast_982_inst_req_1); -- 
    rr_7007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(149), ack => type_cast_982_inst_req_0); -- 
    rr_6984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(149), ack => type_cast_976_inst_req_0); -- 
    cr_6966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(149), ack => type_cast_970_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  place  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	152 
    -- CP-element group 150: 	154 
    -- CP-element group 150: 	156 
    -- CP-element group 150:  members (24) 
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959__entry__
      -- CP-element group 150: 	 branch_block_stmt_223/merge_stmt_917__exit__
      -- CP-element group 150: 	 branch_block_stmt_223/if_stmt_903_else_link/$exit
      -- CP-element group 150: 	 branch_block_stmt_223/if_stmt_903_else_link/else_choice_transition
      -- CP-element group 150: 	 branch_block_stmt_223/ifx_xend_ifx_xelse217
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/$entry
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_update_start_
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_Update/cr
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_update_start_
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_Update/cr
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_update_start_
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_Update/cr
      -- CP-element group 150: 	 branch_block_stmt_223/ifx_xend_ifx_xelse217_PhiReq/$entry
      -- CP-element group 150: 	 branch_block_stmt_223/ifx_xend_ifx_xelse217_PhiReq/$exit
      -- CP-element group 150: 	 branch_block_stmt_223/merge_stmt_917_PhiReqMerge
      -- CP-element group 150: 	 branch_block_stmt_223/merge_stmt_917_PhiAck/$entry
      -- CP-element group 150: 	 branch_block_stmt_223/merge_stmt_917_PhiAck/$exit
      -- CP-element group 150: 	 branch_block_stmt_223/merge_stmt_917_PhiAck/dummy
      -- 
    else_choice_transition_2269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_903_branch_ack_0, ack => zeropad3D_CP_676_elements(150)); -- 
    rr_2285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(150), ack => type_cast_927_inst_req_0); -- 
    cr_2290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(150), ack => type_cast_927_inst_req_1); -- 
    cr_2304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(150), ack => type_cast_936_inst_req_1); -- 
    cr_2318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(150), ack => type_cast_953_inst_req_1); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_Sample/ra
      -- 
    ra_2286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_0, ack => zeropad3D_CP_676_elements(151)); -- 
    -- CP-element group 152:  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (6) 
      -- CP-element group 152: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_927_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_Sample/rr
      -- 
    ca_2291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_1, ack => zeropad3D_CP_676_elements(152)); -- 
    rr_2299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(152), ack => type_cast_936_inst_req_0); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_Sample/ra
      -- 
    ra_2300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_936_inst_ack_0, ack => zeropad3D_CP_676_elements(153)); -- 
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	150 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_936_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_Sample/rr
      -- 
    ca_2305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_936_inst_ack_1, ack => zeropad3D_CP_676_elements(154)); -- 
    rr_2313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(154), ack => type_cast_953_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_Sample/ra
      -- 
    ra_2314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_953_inst_ack_0, ack => zeropad3D_CP_676_elements(155)); -- 
    -- CP-element group 156:  branch  transition  place  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	150 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (13) 
      -- CP-element group 156: 	 branch_block_stmt_223/if_stmt_960__entry__
      -- CP-element group 156: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959__exit__
      -- CP-element group 156: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/$exit
      -- CP-element group 156: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_223/assign_stmt_923_to_assign_stmt_959/type_cast_953_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_223/if_stmt_960_dead_link/$entry
      -- CP-element group 156: 	 branch_block_stmt_223/if_stmt_960_eval_test/$entry
      -- CP-element group 156: 	 branch_block_stmt_223/if_stmt_960_eval_test/$exit
      -- CP-element group 156: 	 branch_block_stmt_223/if_stmt_960_eval_test/branch_req
      -- CP-element group 156: 	 branch_block_stmt_223/R_cmp245_961_place
      -- CP-element group 156: 	 branch_block_stmt_223/if_stmt_960_if_link/$entry
      -- CP-element group 156: 	 branch_block_stmt_223/if_stmt_960_else_link/$entry
      -- 
    ca_2319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_953_inst_ack_1, ack => zeropad3D_CP_676_elements(156)); -- 
    branch_req_2327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(156), ack => if_stmt_960_branch_req_0); -- 
    -- CP-element group 157:  fork  transition  place  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: 	160 
    -- CP-element group 157: 	161 
    -- CP-element group 157: 	162 
    -- CP-element group 157: 	164 
    -- CP-element group 157:  members (33) 
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031__entry__
      -- CP-element group 157: 	 branch_block_stmt_223/merge_stmt_988__exit__
      -- CP-element group 157: 	 branch_block_stmt_223/if_stmt_960_if_link/$exit
      -- CP-element group 157: 	 branch_block_stmt_223/if_stmt_960_if_link/if_choice_transition
      -- CP-element group 157: 	 branch_block_stmt_223/ifx_xelse217_whilex_xend
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_update_start_
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_Sample/rr
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_update_start_
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_word_address_calculated
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_root_address_calculated
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Sample/word_access_start/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Sample/word_access_start/word_0/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Sample/word_access_start/word_0/rr
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/word_access_complete/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/word_access_complete/word_0/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/word_access_complete/word_0/cr
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_update_start_
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_223/merge_stmt_988_PhiAck/dummy
      -- CP-element group 157: 	 branch_block_stmt_223/merge_stmt_988_PhiAck/$exit
      -- CP-element group 157: 	 branch_block_stmt_223/merge_stmt_988_PhiAck/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/ifx_xelse217_whilex_xend_PhiReq/$exit
      -- CP-element group 157: 	 branch_block_stmt_223/ifx_xelse217_whilex_xend_PhiReq/$entry
      -- CP-element group 157: 	 branch_block_stmt_223/merge_stmt_988_PhiReqMerge
      -- 
    if_choice_transition_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_960_branch_ack_1, ack => zeropad3D_CP_676_elements(157)); -- 
    rr_2349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(157), ack => type_cast_991_inst_req_0); -- 
    cr_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(157), ack => type_cast_991_inst_req_1); -- 
    rr_2371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(157), ack => LOAD_pad_1000_load_0_req_0); -- 
    cr_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(157), ack => LOAD_pad_1000_load_0_req_1); -- 
    cr_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(157), ack => type_cast_1004_inst_req_1); -- 
    -- CP-element group 158:  fork  transition  place  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	606 
    -- CP-element group 158: 	607 
    -- CP-element group 158: 	609 
    -- CP-element group 158: 	610 
    -- CP-element group 158: 	612 
    -- CP-element group 158:  members (22) 
      -- CP-element group 158: 	 branch_block_stmt_223/if_stmt_960_else_link/$exit
      -- CP-element group 158: 	 branch_block_stmt_223/if_stmt_960_else_link/else_choice_transition
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/SplitProtocol/Update/cr
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/SplitProtocol/Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/SplitProtocol/Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_979/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/SplitProtocol/Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/SplitProtocol/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/SplitProtocol/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/SplitProtocol/Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/SplitProtocol/Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/SplitProtocol/Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/SplitProtocol/Update/cr
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/$entry
      -- CP-element group 158: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/$entry
      -- 
    else_choice_transition_2336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_960_branch_ack_0, ack => zeropad3D_CP_676_elements(158)); -- 
    cr_6932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(158), ack => type_cast_978_inst_req_1); -- 
    rr_6927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(158), ack => type_cast_978_inst_req_0); -- 
    rr_6904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(158), ack => type_cast_972_inst_req_0); -- 
    cr_6909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(158), ack => type_cast_972_inst_req_1); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_Sample/ra
      -- 
    ra_2350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_991_inst_ack_0, ack => zeropad3D_CP_676_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	157 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	165 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_991_Update/ca
      -- 
    ca_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_991_inst_ack_1, ack => zeropad3D_CP_676_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	157 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (5) 
      -- CP-element group 161: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Sample/word_access_start/$exit
      -- CP-element group 161: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Sample/word_access_start/word_0/$exit
      -- CP-element group 161: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Sample/word_access_start/word_0/ra
      -- 
    ra_2372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1000_load_0_ack_0, ack => zeropad3D_CP_676_elements(161)); -- 
    -- CP-element group 162:  transition  input  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	157 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (12) 
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/word_access_complete/$exit
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/word_access_complete/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/word_access_complete/word_0/ca
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/LOAD_pad_1000_Merge/$entry
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/LOAD_pad_1000_Merge/$exit
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/LOAD_pad_1000_Merge/merge_req
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/LOAD_pad_1000_Update/LOAD_pad_1000_Merge/merge_ack
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_Sample/rr
      -- 
    ca_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1000_load_0_ack_1, ack => zeropad3D_CP_676_elements(162)); -- 
    rr_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(162), ack => type_cast_1004_inst_req_0); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_Sample/ra
      -- 
    ra_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1004_inst_ack_0, ack => zeropad3D_CP_676_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	157 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/type_cast_1004_Update/ca
      -- 
    ca_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1004_inst_ack_1, ack => zeropad3D_CP_676_elements(164)); -- 
    -- CP-element group 165:  join  fork  transition  place  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	160 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	639 
    -- CP-element group 165: 	640 
    -- CP-element group 165: 	642 
    -- CP-element group 165: 	643 
    -- CP-element group 165:  members (16) 
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313
      -- CP-element group 165: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031__exit__
      -- CP-element group 165: 	 branch_block_stmt_223/assign_stmt_992_to_assign_stmt_1031/$exit
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/SplitProtocol/Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/SplitProtocol/Sample/rr
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/SplitProtocol/$entry
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/$entry
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/$entry
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/$entry
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/$entry
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/$entry
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1047/$entry
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1040/$entry
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/SplitProtocol/Update/cr
      -- CP-element group 165: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/SplitProtocol/Update/$entry
      -- 
    rr_7120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(165), ack => type_cast_1037_inst_req_0); -- 
    cr_7125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(165), ack => type_cast_1037_inst_req_1); -- 
    zeropad3D_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(160) & zeropad3D_CP_676_elements(164);
      gj_zeropad3D_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	649 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_Sample/ra
      -- 
    ra_2414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1058_inst_ack_0, ack => zeropad3D_CP_676_elements(166)); -- 
    -- CP-element group 167:  branch  transition  place  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	649 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (13) 
      -- CP-element group 167: 	 branch_block_stmt_223/if_stmt_1085__entry__
      -- CP-element group 167: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084__exit__
      -- CP-element group 167: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/$exit
      -- CP-element group 167: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_Update/ca
      -- CP-element group 167: 	 branch_block_stmt_223/if_stmt_1085_dead_link/$entry
      -- CP-element group 167: 	 branch_block_stmt_223/if_stmt_1085_eval_test/$entry
      -- CP-element group 167: 	 branch_block_stmt_223/if_stmt_1085_eval_test/$exit
      -- CP-element group 167: 	 branch_block_stmt_223/if_stmt_1085_eval_test/branch_req
      -- CP-element group 167: 	 branch_block_stmt_223/R_orx_xcond1850_1086_place
      -- CP-element group 167: 	 branch_block_stmt_223/if_stmt_1085_if_link/$entry
      -- CP-element group 167: 	 branch_block_stmt_223/if_stmt_1085_else_link/$entry
      -- 
    ca_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1058_inst_ack_1, ack => zeropad3D_CP_676_elements(167)); -- 
    branch_req_2427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => if_stmt_1085_branch_req_0); -- 
    -- CP-element group 168:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: 	171 
    -- CP-element group 168:  members (18) 
      -- CP-element group 168: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121__entry__
      -- CP-element group 168: 	 branch_block_stmt_223/merge_stmt_1091__exit__
      -- CP-element group 168: 	 branch_block_stmt_223/if_stmt_1085_if_link/$exit
      -- CP-element group 168: 	 branch_block_stmt_223/if_stmt_1085_if_link/if_choice_transition
      -- CP-element group 168: 	 branch_block_stmt_223/whilex_xbody313_lorx_xlhsx_xfalse331
      -- CP-element group 168: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/$entry
      -- CP-element group 168: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_update_start_
      -- CP-element group 168: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_Sample/rr
      -- CP-element group 168: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_Update/cr
      -- CP-element group 168: 	 branch_block_stmt_223/merge_stmt_1091_PhiAck/$entry
      -- CP-element group 168: 	 branch_block_stmt_223/whilex_xbody313_lorx_xlhsx_xfalse331_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_223/merge_stmt_1091_PhiAck/dummy
      -- CP-element group 168: 	 branch_block_stmt_223/merge_stmt_1091_PhiAck/$exit
      -- CP-element group 168: 	 branch_block_stmt_223/whilex_xbody313_lorx_xlhsx_xfalse331_PhiReq/$exit
      -- CP-element group 168: 	 branch_block_stmt_223/merge_stmt_1091_PhiReqMerge
      -- 
    if_choice_transition_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1085_branch_ack_1, ack => zeropad3D_CP_676_elements(168)); -- 
    rr_2449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(168), ack => type_cast_1095_inst_req_0); -- 
    cr_2454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(168), ack => type_cast_1095_inst_req_1); -- 
    -- CP-element group 169:  transition  place  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	650 
    -- CP-element group 169:  members (5) 
      -- CP-element group 169: 	 branch_block_stmt_223/if_stmt_1085_else_link/$exit
      -- CP-element group 169: 	 branch_block_stmt_223/if_stmt_1085_else_link/else_choice_transition
      -- CP-element group 169: 	 branch_block_stmt_223/whilex_xbody313_ifx_xthen348
      -- CP-element group 169: 	 branch_block_stmt_223/whilex_xbody313_ifx_xthen348_PhiReq/$exit
      -- CP-element group 169: 	 branch_block_stmt_223/whilex_xbody313_ifx_xthen348_PhiReq/$entry
      -- 
    else_choice_transition_2436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1085_branch_ack_0, ack => zeropad3D_CP_676_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_Sample/ra
      -- 
    ra_2450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1095_inst_ack_0, ack => zeropad3D_CP_676_elements(170)); -- 
    -- CP-element group 171:  branch  transition  place  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	168 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (13) 
      -- CP-element group 171: 	 branch_block_stmt_223/if_stmt_1122__entry__
      -- CP-element group 171: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121__exit__
      -- CP-element group 171: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/$exit
      -- CP-element group 171: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_223/assign_stmt_1096_to_assign_stmt_1121/type_cast_1095_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_223/if_stmt_1122_dead_link/$entry
      -- CP-element group 171: 	 branch_block_stmt_223/if_stmt_1122_eval_test/$entry
      -- CP-element group 171: 	 branch_block_stmt_223/if_stmt_1122_eval_test/$exit
      -- CP-element group 171: 	 branch_block_stmt_223/if_stmt_1122_eval_test/branch_req
      -- CP-element group 171: 	 branch_block_stmt_223/R_orx_xcond1851_1123_place
      -- CP-element group 171: 	 branch_block_stmt_223/if_stmt_1122_if_link/$entry
      -- CP-element group 171: 	 branch_block_stmt_223/if_stmt_1122_else_link/$entry
      -- 
    ca_2455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1095_inst_ack_1, ack => zeropad3D_CP_676_elements(171)); -- 
    branch_req_2463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(171), ack => if_stmt_1122_branch_req_0); -- 
    -- CP-element group 172:  fork  transition  place  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	188 
    -- CP-element group 172: 	189 
    -- CP-element group 172: 	191 
    -- CP-element group 172: 	193 
    -- CP-element group 172: 	195 
    -- CP-element group 172: 	197 
    -- CP-element group 172: 	199 
    -- CP-element group 172: 	201 
    -- CP-element group 172: 	203 
    -- CP-element group 172: 	206 
    -- CP-element group 172:  members (46) 
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Update/word_access_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_complete/req
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291__entry__
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/merge_stmt_1186__exit__
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/word_access_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_update_start_
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_complete/req
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_final_index_sum_regn_update_start
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/word_access_complete/word_0/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_complete/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Update/word_access_complete/word_0/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_final_index_sum_regn_Update/req
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_final_index_sum_regn_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_final_index_sum_regn_update_start
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_final_index_sum_regn_Update/req
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_update_start_
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_final_index_sum_regn_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_update_start_
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_update_start_
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Update/word_access_complete/word_0/cr
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/word_access_complete/word_0/cr
      -- CP-element group 172: 	 branch_block_stmt_223/if_stmt_1122_if_link/$exit
      -- CP-element group 172: 	 branch_block_stmt_223/if_stmt_1122_if_link/if_choice_transition
      -- CP-element group 172: 	 branch_block_stmt_223/lorx_xlhsx_xfalse331_ifx_xelse369
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_update_start_
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_update_start_
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_update_start_
      -- CP-element group 172: 	 branch_block_stmt_223/merge_stmt_1186_PhiAck/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/merge_stmt_1186_PhiAck/$exit
      -- CP-element group 172: 	 branch_block_stmt_223/lorx_xlhsx_xfalse331_ifx_xelse369_PhiReq/$exit
      -- CP-element group 172: 	 branch_block_stmt_223/lorx_xlhsx_xfalse331_ifx_xelse369_PhiReq/$entry
      -- CP-element group 172: 	 branch_block_stmt_223/merge_stmt_1186_PhiReqMerge
      -- CP-element group 172: 	 branch_block_stmt_223/merge_stmt_1186_PhiAck/dummy
      -- 
    if_choice_transition_2468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1122_branch_ack_1, ack => zeropad3D_CP_676_elements(172)); -- 
    req_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => addr_of_1286_final_reg_req_1); -- 
    req_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => addr_of_1261_final_reg_req_1); -- 
    req_2786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => array_obj_ref_1285_index_offset_req_1); -- 
    req_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => array_obj_ref_1260_index_offset_req_1); -- 
    cr_2755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => type_cast_1279_inst_req_1); -- 
    cr_2851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => ptr_deref_1289_store_0_req_1); -- 
    cr_2736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => ptr_deref_1265_load_0_req_1); -- 
    rr_2626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => type_cast_1190_inst_req_0); -- 
    cr_2631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => type_cast_1190_inst_req_1); -- 
    cr_2645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(172), ack => type_cast_1254_inst_req_1); -- 
    -- CP-element group 173:  transition  place  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	650 
    -- CP-element group 173:  members (5) 
      -- CP-element group 173: 	 branch_block_stmt_223/if_stmt_1122_else_link/$exit
      -- CP-element group 173: 	 branch_block_stmt_223/if_stmt_1122_else_link/else_choice_transition
      -- CP-element group 173: 	 branch_block_stmt_223/lorx_xlhsx_xfalse331_ifx_xthen348
      -- CP-element group 173: 	 branch_block_stmt_223/lorx_xlhsx_xfalse331_ifx_xthen348_PhiReq/$exit
      -- CP-element group 173: 	 branch_block_stmt_223/lorx_xlhsx_xfalse331_ifx_xthen348_PhiReq/$entry
      -- 
    else_choice_transition_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1122_branch_ack_0, ack => zeropad3D_CP_676_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	650 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_Sample/ra
      -- 
    ra_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1132_inst_ack_0, ack => zeropad3D_CP_676_elements(174)); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	650 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	178 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_Update/ca
      -- 
    ca_2491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1132_inst_ack_1, ack => zeropad3D_CP_676_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	650 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_Sample/ra
      -- 
    ra_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1137_inst_ack_0, ack => zeropad3D_CP_676_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	650 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_Update/ca
      -- 
    ca_2505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1137_inst_ack_1, ack => zeropad3D_CP_676_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	175 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_Sample/rr
      -- 
    rr_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(178), ack => type_cast_1171_inst_req_0); -- 
    zeropad3D_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(175) & zeropad3D_CP_676_elements(177);
      gj_zeropad3D_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_Sample/ra
      -- 
    ra_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_0, ack => zeropad3D_CP_676_elements(179)); -- 
    -- CP-element group 180:  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	650 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (16) 
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_resized_1
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_scaled_1
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_computed_1
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_resize_1/$entry
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_resize_1/$exit
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_resize_1/index_resize_req
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_resize_1/index_resize_ack
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_scale_1/$entry
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_scale_1/$exit
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_scale_1/scale_rename_req
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_index_scale_1/scale_rename_ack
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_final_index_sum_regn_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_final_index_sum_regn_Sample/req
      -- 
    ca_2519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_1, ack => zeropad3D_CP_676_elements(180)); -- 
    req_2544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(180), ack => array_obj_ref_1177_index_offset_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	187 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_final_index_sum_regn_sample_complete
      -- CP-element group 181: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_final_index_sum_regn_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_final_index_sum_regn_Sample/ack
      -- 
    ack_2545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1177_index_offset_ack_0, ack => zeropad3D_CP_676_elements(181)); -- 
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	650 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (11) 
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_root_address_calculated
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_offset_calculated
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_final_index_sum_regn_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_final_index_sum_regn_Update/ack
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_base_plus_offset/$entry
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_base_plus_offset/$exit
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_base_plus_offset/sum_rename_req
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_base_plus_offset/sum_rename_ack
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_request/$entry
      -- CP-element group 182: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_request/req
      -- 
    ack_2550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1177_index_offset_ack_1, ack => zeropad3D_CP_676_elements(182)); -- 
    req_2559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(182), ack => addr_of_1178_final_reg_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_request/$exit
      -- CP-element group 183: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_request/ack
      -- 
    ack_2560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1178_final_reg_ack_0, ack => zeropad3D_CP_676_elements(183)); -- 
    -- CP-element group 184:  join  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	650 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (28) 
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_complete/$exit
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_complete/ack
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_base_address_calculated
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_word_address_calculated
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_root_address_calculated
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_base_address_resized
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_base_addr_resize/$entry
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_base_addr_resize/$exit
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_base_addr_resize/base_resize_req
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_base_addr_resize/base_resize_ack
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_base_plus_offset/$entry
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_base_plus_offset/$exit
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_base_plus_offset/sum_rename_req
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_base_plus_offset/sum_rename_ack
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_word_addrgen/$entry
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_word_addrgen/$exit
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_word_addrgen/root_register_req
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_word_addrgen/root_register_ack
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/ptr_deref_1181_Split/$entry
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/ptr_deref_1181_Split/$exit
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/ptr_deref_1181_Split/split_req
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/ptr_deref_1181_Split/split_ack
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/word_access_start/$entry
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/word_access_start/word_0/$entry
      -- CP-element group 184: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/word_access_start/word_0/rr
      -- 
    ack_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1178_final_reg_ack_1, ack => zeropad3D_CP_676_elements(184)); -- 
    rr_2603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(184), ack => ptr_deref_1181_store_0_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (5) 
      -- CP-element group 185: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/word_access_start/$exit
      -- CP-element group 185: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/word_access_start/word_0/$exit
      -- CP-element group 185: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Sample/word_access_start/word_0/ra
      -- 
    ra_2604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1181_store_0_ack_0, ack => zeropad3D_CP_676_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	650 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (5) 
      -- CP-element group 186: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Update/word_access_complete/$exit
      -- CP-element group 186: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Update/word_access_complete/word_0/$exit
      -- CP-element group 186: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Update/word_access_complete/word_0/ca
      -- 
    ca_2615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1181_store_0_ack_1, ack => zeropad3D_CP_676_elements(186)); -- 
    -- CP-element group 187:  join  transition  place  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	181 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	651 
    -- CP-element group 187:  members (5) 
      -- CP-element group 187: 	 branch_block_stmt_223/ifx_xthen348_ifx_xend417
      -- CP-element group 187: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184__exit__
      -- CP-element group 187: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/$exit
      -- CP-element group 187: 	 branch_block_stmt_223/ifx_xthen348_ifx_xend417_PhiReq/$exit
      -- CP-element group 187: 	 branch_block_stmt_223/ifx_xthen348_ifx_xend417_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(181) & zeropad3D_CP_676_elements(186);
      gj_zeropad3D_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	172 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_Sample/ra
      -- 
    ra_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1190_inst_ack_0, ack => zeropad3D_CP_676_elements(188)); -- 
    -- CP-element group 189:  fork  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	172 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189: 	198 
    -- CP-element group 189:  members (9) 
      -- CP-element group 189: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_Sample/rr
      -- CP-element group 189: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1190_Update/ca
      -- CP-element group 189: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_Sample/rr
      -- 
    ca_2632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1190_inst_ack_1, ack => zeropad3D_CP_676_elements(189)); -- 
    rr_2640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(189), ack => type_cast_1254_inst_req_0); -- 
    rr_2750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(189), ack => type_cast_1279_inst_req_0); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_Sample/ra
      -- 
    ra_2641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1254_inst_ack_0, ack => zeropad3D_CP_676_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	172 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (16) 
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_final_index_sum_regn_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_scale_1/scale_rename_req
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_scale_1/$entry
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_scale_1/$exit
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_scale_1/scale_rename_ack
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_resize_1/index_resize_ack
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_resize_1/index_resize_req
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_resize_1/$exit
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_resize_1/$entry
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_computed_1
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_final_index_sum_regn_Sample/req
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_scaled_1
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_index_resized_1
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1254_Update/ca
      -- 
    ca_2646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1254_inst_ack_1, ack => zeropad3D_CP_676_elements(191)); -- 
    req_2671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(191), ack => array_obj_ref_1260_index_offset_req_0); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	207 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_final_index_sum_regn_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_final_index_sum_regn_sample_complete
      -- CP-element group 192: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_final_index_sum_regn_Sample/ack
      -- 
    ack_2672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1260_index_offset_ack_0, ack => zeropad3D_CP_676_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	172 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (11) 
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_request/req
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_request/$entry
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_base_plus_offset/sum_rename_ack
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_base_plus_offset/sum_rename_req
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_base_plus_offset/$exit
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_base_plus_offset/$entry
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_final_index_sum_regn_Update/ack
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_final_index_sum_regn_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_offset_calculated
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1260_root_address_calculated
      -- 
    ack_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1260_index_offset_ack_1, ack => zeropad3D_CP_676_elements(193)); -- 
    req_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(193), ack => addr_of_1261_final_reg_req_0); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_request/ack
      -- CP-element group 194: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_request/$exit
      -- CP-element group 194: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_sample_completed_
      -- 
    ack_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1261_final_reg_ack_0, ack => zeropad3D_CP_676_elements(194)); -- 
    -- CP-element group 195:  join  fork  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	172 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (24) 
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_complete/$exit
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_base_plus_offset/sum_rename_req
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_word_addrgen/$exit
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_base_plus_offset/sum_rename_ack
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_word_addrgen/root_register_req
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_word_addrgen/root_register_ack
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_word_addrgen/$entry
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_base_plus_offset/$exit
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_base_plus_offset/$entry
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_base_addr_resize/base_resize_ack
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_base_addr_resize/$exit
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Sample/word_access_start/word_0/rr
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_base_addr_resize/base_resize_req
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Sample/word_access_start/word_0/$entry
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_base_addr_resize/$entry
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Sample/word_access_start/$entry
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_base_address_resized
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_root_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_word_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_base_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_complete/ack
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1261_update_completed_
      -- 
    ack_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1261_final_reg_ack_1, ack => zeropad3D_CP_676_elements(195)); -- 
    rr_2725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(195), ack => ptr_deref_1265_load_0_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (5) 
      -- CP-element group 196: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Sample/word_access_start/word_0/ra
      -- CP-element group 196: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Sample/word_access_start/word_0/$exit
      -- CP-element group 196: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Sample/word_access_start/$exit
      -- CP-element group 196: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Sample/$exit
      -- 
    ra_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1265_load_0_ack_0, ack => zeropad3D_CP_676_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	172 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	204 
    -- CP-element group 197:  members (9) 
      -- CP-element group 197: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/word_access_complete/$exit
      -- CP-element group 197: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/word_access_complete/word_0/$exit
      -- CP-element group 197: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/ptr_deref_1265_Merge/merge_ack
      -- CP-element group 197: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/ptr_deref_1265_Merge/merge_req
      -- CP-element group 197: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/ptr_deref_1265_Merge/$exit
      -- CP-element group 197: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/ptr_deref_1265_Merge/$entry
      -- CP-element group 197: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1265_Update/word_access_complete/word_0/ca
      -- 
    ca_2737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1265_load_0_ack_1, ack => zeropad3D_CP_676_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	189 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_sample_completed_
      -- 
    ra_2751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_0, ack => zeropad3D_CP_676_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	172 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (16) 
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_final_index_sum_regn_Sample/req
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_final_index_sum_regn_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_scale_1/scale_rename_ack
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_scale_1/scale_rename_req
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_scale_1/$exit
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_scale_1/$entry
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_resize_1/index_resize_ack
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_resize_1/index_resize_req
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_resize_1/$exit
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_resize_1/$entry
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_computed_1
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_scaled_1
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_index_resized_1
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_Update/ca
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/type_cast_1279_update_completed_
      -- 
    ca_2756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_1, ack => zeropad3D_CP_676_elements(199)); -- 
    req_2781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(199), ack => array_obj_ref_1285_index_offset_req_0); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	207 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_final_index_sum_regn_Sample/ack
      -- CP-element group 200: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_final_index_sum_regn_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_final_index_sum_regn_sample_complete
      -- 
    ack_2782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1285_index_offset_ack_0, ack => zeropad3D_CP_676_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	172 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (11) 
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_request/req
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_base_plus_offset/$exit
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_base_plus_offset/sum_rename_req
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_final_index_sum_regn_Update/ack
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_base_plus_offset/sum_rename_ack
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_base_plus_offset/$entry
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_request/$entry
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_final_index_sum_regn_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_offset_calculated
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/array_obj_ref_1285_root_address_calculated
      -- CP-element group 201: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_sample_start_
      -- 
    ack_2787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1285_index_offset_ack_1, ack => zeropad3D_CP_676_elements(201)); -- 
    req_2796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(201), ack => addr_of_1286_final_reg_req_0); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_request/ack
      -- CP-element group 202: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_request/$exit
      -- CP-element group 202: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_sample_completed_
      -- 
    ack_2797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1286_final_reg_ack_0, ack => zeropad3D_CP_676_elements(202)); -- 
    -- CP-element group 203:  fork  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	172 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (19) 
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_base_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_complete/$exit
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_complete/ack
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_word_addrgen/root_register_ack
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/addr_of_1286_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_word_addrgen/root_register_req
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_word_addrgen/$exit
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_word_addrgen/$entry
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_base_plus_offset/sum_rename_ack
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_base_plus_offset/sum_rename_req
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_base_plus_offset/$exit
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_base_plus_offset/$entry
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_base_addr_resize/base_resize_ack
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_base_addr_resize/base_resize_req
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_base_addr_resize/$exit
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_base_addr_resize/$entry
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_base_address_resized
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_root_address_calculated
      -- CP-element group 203: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_word_address_calculated
      -- 
    ack_2802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1286_final_reg_ack_1, ack => zeropad3D_CP_676_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	197 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (9) 
      -- CP-element group 204: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/word_access_start/word_0/rr
      -- CP-element group 204: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/word_access_start/word_0/$entry
      -- CP-element group 204: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/word_access_start/$entry
      -- CP-element group 204: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/ptr_deref_1289_Split/split_ack
      -- CP-element group 204: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/ptr_deref_1289_Split/split_req
      -- CP-element group 204: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/ptr_deref_1289_Split/$exit
      -- CP-element group 204: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/ptr_deref_1289_Split/$entry
      -- CP-element group 204: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/$entry
      -- 
    rr_2840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(204), ack => ptr_deref_1289_store_0_req_0); -- 
    zeropad3D_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(197) & zeropad3D_CP_676_elements(203);
      gj_zeropad3D_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (5) 
      -- CP-element group 205: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/word_access_start/word_0/$exit
      -- CP-element group 205: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/word_access_start/word_0/ra
      -- CP-element group 205: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/word_access_start/$exit
      -- CP-element group 205: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Sample/$exit
      -- 
    ra_2841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1289_store_0_ack_0, ack => zeropad3D_CP_676_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	172 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Update/word_access_complete/$exit
      -- CP-element group 206: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Update/word_access_complete/word_0/ca
      -- CP-element group 206: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/ptr_deref_1289_Update/word_access_complete/word_0/$exit
      -- 
    ca_2852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1289_store_0_ack_1, ack => zeropad3D_CP_676_elements(206)); -- 
    -- CP-element group 207:  join  transition  place  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	192 
    -- CP-element group 207: 	200 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	651 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_223/ifx_xelse369_ifx_xend417
      -- CP-element group 207: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291__exit__
      -- CP-element group 207: 	 branch_block_stmt_223/assign_stmt_1191_to_assign_stmt_1291/$exit
      -- CP-element group 207: 	 branch_block_stmt_223/ifx_xelse369_ifx_xend417_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_223/ifx_xelse369_ifx_xend417_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(192) & zeropad3D_CP_676_elements(200) & zeropad3D_CP_676_elements(206);
      gj_zeropad3D_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	651 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_Sample/ra
      -- CP-element group 208: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_sample_completed_
      -- 
    ra_2864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1297_inst_ack_0, ack => zeropad3D_CP_676_elements(208)); -- 
    -- CP-element group 209:  branch  transition  place  input  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	651 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311__exit__
      -- CP-element group 209: 	 branch_block_stmt_223/if_stmt_1312__entry__
      -- CP-element group 209: 	 branch_block_stmt_223/if_stmt_1312_else_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_223/if_stmt_1312_if_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_223/if_stmt_1312_eval_test/branch_req
      -- CP-element group 209: 	 branch_block_stmt_223/if_stmt_1312_eval_test/$exit
      -- CP-element group 209: 	 branch_block_stmt_223/if_stmt_1312_eval_test/$entry
      -- CP-element group 209: 	 branch_block_stmt_223/if_stmt_1312_dead_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_Update/ca
      -- CP-element group 209: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/$exit
      -- CP-element group 209: 	 branch_block_stmt_223/R_cmp425_1313_place
      -- 
    ca_2869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1297_inst_ack_1, ack => zeropad3D_CP_676_elements(209)); -- 
    branch_req_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(209), ack => if_stmt_1312_branch_req_0); -- 
    -- CP-element group 210:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	660 
    -- CP-element group 210: 	661 
    -- CP-element group 210: 	663 
    -- CP-element group 210: 	664 
    -- CP-element group 210: 	666 
    -- CP-element group 210: 	667 
    -- CP-element group 210:  members (40) 
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468
      -- CP-element group 210: 	 branch_block_stmt_223/assign_stmt_1324__exit__
      -- CP-element group 210: 	 branch_block_stmt_223/assign_stmt_1324__entry__
      -- CP-element group 210: 	 branch_block_stmt_223/merge_stmt_1318__exit__
      -- CP-element group 210: 	 branch_block_stmt_223/assign_stmt_1324/$exit
      -- CP-element group 210: 	 branch_block_stmt_223/assign_stmt_1324/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/if_stmt_1312_if_link/if_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_223/if_stmt_1312_if_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xend417_ifx_xthen427
      -- CP-element group 210: 	 branch_block_stmt_223/merge_stmt_1318_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/merge_stmt_1318_PhiAck/dummy
      -- CP-element group 210: 	 branch_block_stmt_223/merge_stmt_1318_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_223/merge_stmt_1318_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xend417_ifx_xthen427_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xend417_ifx_xthen427_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/SplitProtocol/Update/cr
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/SplitProtocol/Update/cr
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1312_branch_ack_1, ack => zeropad3D_CP_676_elements(210)); -- 
    rr_7296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(210), ack => type_cast_1378_inst_req_0); -- 
    cr_7301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(210), ack => type_cast_1378_inst_req_1); -- 
    rr_7319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(210), ack => type_cast_1384_inst_req_0); -- 
    cr_7324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(210), ack => type_cast_1384_inst_req_1); -- 
    rr_7342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(210), ack => type_cast_1390_inst_req_0); -- 
    cr_7347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(210), ack => type_cast_1390_inst_req_1); -- 
    -- CP-element group 211:  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211: 	213 
    -- CP-element group 211: 	215 
    -- CP-element group 211: 	217 
    -- CP-element group 211:  members (24) 
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367__entry__
      -- CP-element group 211: 	 branch_block_stmt_223/merge_stmt_1326__exit__
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_update_start_
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_Update/cr
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_Update/cr
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_update_start_
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/$entry
      -- CP-element group 211: 	 branch_block_stmt_223/if_stmt_1312_else_link/else_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_223/if_stmt_1312_else_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_Update/cr
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_update_start_
      -- CP-element group 211: 	 branch_block_stmt_223/ifx_xend417_ifx_xelse432
      -- CP-element group 211: 	 branch_block_stmt_223/merge_stmt_1326_PhiReqMerge
      -- CP-element group 211: 	 branch_block_stmt_223/merge_stmt_1326_PhiAck/dummy
      -- CP-element group 211: 	 branch_block_stmt_223/merge_stmt_1326_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_223/merge_stmt_1326_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_223/ifx_xend417_ifx_xelse432_PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_223/ifx_xend417_ifx_xelse432_PhiReq/$entry
      -- 
    else_choice_transition_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1312_branch_ack_0, ack => zeropad3D_CP_676_elements(211)); -- 
    cr_2921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(211), ack => type_cast_1345_inst_req_1); -- 
    cr_2907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(211), ack => type_cast_1336_inst_req_1); -- 
    rr_2902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(211), ack => type_cast_1336_inst_req_0); -- 
    cr_2935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(211), ack => type_cast_1361_inst_req_1); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_Sample/ra
      -- CP-element group 212: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_sample_completed_
      -- 
    ra_2903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1336_inst_ack_0, ack => zeropad3D_CP_676_elements(212)); -- 
    -- CP-element group 213:  transition  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (6) 
      -- CP-element group 213: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_Sample/rr
      -- CP-element group 213: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_sample_start_
      -- CP-element group 213: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_Sample/$entry
      -- CP-element group 213: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_Update/ca
      -- CP-element group 213: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1336_update_completed_
      -- 
    ca_2908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1336_inst_ack_1, ack => zeropad3D_CP_676_elements(213)); -- 
    rr_2916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(213), ack => type_cast_1345_inst_req_0); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_sample_completed_
      -- CP-element group 214: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_Sample/ra
      -- CP-element group 214: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_Sample/$exit
      -- 
    ra_2917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1345_inst_ack_0, ack => zeropad3D_CP_676_elements(214)); -- 
    -- CP-element group 215:  transition  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	211 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_Update/$exit
      -- CP-element group 215: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1345_Update/ca
      -- CP-element group 215: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_Sample/rr
      -- CP-element group 215: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_sample_start_
      -- 
    ca_2922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1345_inst_ack_1, ack => zeropad3D_CP_676_elements(215)); -- 
    rr_2930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(215), ack => type_cast_1361_inst_req_0); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_Sample/ra
      -- CP-element group 216: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_sample_completed_
      -- 
    ra_2931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_0, ack => zeropad3D_CP_676_elements(216)); -- 
    -- CP-element group 217:  branch  transition  place  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	211 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (13) 
      -- CP-element group 217: 	 branch_block_stmt_223/if_stmt_1368__entry__
      -- CP-element group 217: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367__exit__
      -- CP-element group 217: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/$exit
      -- CP-element group 217: 	 branch_block_stmt_223/if_stmt_1368_else_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_223/if_stmt_1368_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_223/if_stmt_1368_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_223/if_stmt_1368_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_223/if_stmt_1368_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_223/if_stmt_1368_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_Update/ca
      -- CP-element group 217: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_223/R_cmp459_1369_place
      -- CP-element group 217: 	 branch_block_stmt_223/assign_stmt_1332_to_assign_stmt_1367/type_cast_1361_update_completed_
      -- 
    ca_2936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_1, ack => zeropad3D_CP_676_elements(217)); -- 
    branch_req_2944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(217), ack => if_stmt_1368_branch_req_0); -- 
    -- CP-element group 218:  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218: 	222 
    -- CP-element group 218: 	223 
    -- CP-element group 218: 	225 
    -- CP-element group 218:  members (33) 
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Sample/word_access_start/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445__entry__
      -- CP-element group 218: 	 branch_block_stmt_223/merge_stmt_1396__exit__
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/word_access_complete/word_0/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/word_access_complete/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_root_address_calculated
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_word_address_calculated
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Sample/word_access_start/word_0/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/word_access_complete/word_0/cr
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_update_start_
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_update_start_
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_update_start_
      -- CP-element group 218: 	 branch_block_stmt_223/if_stmt_1368_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_223/if_stmt_1368_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/ifx_xelse432_whilex_xend469
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Sample/word_access_start/word_0/rr
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/merge_stmt_1396_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_223/ifx_xelse432_whilex_xend469_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/ifx_xelse432_whilex_xend469_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_223/merge_stmt_1396_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_223/merge_stmt_1396_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_223/merge_stmt_1396_PhiAck/dummy
      -- 
    if_choice_transition_2949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1368_branch_ack_1, ack => zeropad3D_CP_676_elements(218)); -- 
    cr_2999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(218), ack => LOAD_pad_1408_load_0_req_1); -- 
    cr_2971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(218), ack => type_cast_1399_inst_req_1); -- 
    rr_2966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(218), ack => type_cast_1399_inst_req_0); -- 
    rr_2988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(218), ack => LOAD_pad_1408_load_0_req_0); -- 
    cr_3018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(218), ack => type_cast_1412_inst_req_1); -- 
    -- CP-element group 219:  fork  transition  place  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	652 
    -- CP-element group 219: 	653 
    -- CP-element group 219: 	655 
    -- CP-element group 219: 	656 
    -- CP-element group 219: 	658 
    -- CP-element group 219:  members (22) 
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468
      -- CP-element group 219: 	 branch_block_stmt_223/if_stmt_1368_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_223/if_stmt_1368_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/SplitProtocol/Sample/rr
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/SplitProtocol/Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/SplitProtocol/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/SplitProtocol/Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/SplitProtocol/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1387/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/SplitProtocol/Update/cr
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/SplitProtocol/Update/cr
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/SplitProtocol/Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/SplitProtocol/Sample/rr
      -- CP-element group 219: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/SplitProtocol/Sample/$entry
      -- 
    else_choice_transition_2953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1368_branch_ack_0, ack => zeropad3D_CP_676_elements(219)); -- 
    rr_7239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(219), ack => type_cast_1380_inst_req_0); -- 
    cr_7267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(219), ack => type_cast_1386_inst_req_1); -- 
    cr_7244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(219), ack => type_cast_1380_inst_req_1); -- 
    rr_7262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(219), ack => type_cast_1386_inst_req_0); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_Sample/ra
      -- CP-element group 220: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_sample_completed_
      -- 
    ra_2967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1399_inst_ack_0, ack => zeropad3D_CP_676_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	226 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1399_update_completed_
      -- 
    ca_2972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1399_inst_ack_1, ack => zeropad3D_CP_676_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	218 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (5) 
      -- CP-element group 222: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Sample/word_access_start/$exit
      -- CP-element group 222: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Sample/word_access_start/word_0/$exit
      -- CP-element group 222: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_sample_completed_
      -- CP-element group 222: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Sample/word_access_start/word_0/ra
      -- 
    ra_2989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1408_load_0_ack_0, ack => zeropad3D_CP_676_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	218 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (12) 
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/word_access_complete/word_0/$exit
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_Sample/rr
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/word_access_complete/$exit
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/word_access_complete/word_0/ca
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_Sample/$entry
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/LOAD_pad_1408_Merge/$entry
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/LOAD_pad_1408_Merge/$exit
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_update_completed_
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/LOAD_pad_1408_Merge/merge_ack
      -- CP-element group 223: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/LOAD_pad_1408_Update/LOAD_pad_1408_Merge/merge_req
      -- 
    ca_3000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1408_load_0_ack_1, ack => zeropad3D_CP_676_elements(223)); -- 
    rr_3013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(223), ack => type_cast_1412_inst_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_Sample/ra
      -- 
    ra_3014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1412_inst_ack_0, ack => zeropad3D_CP_676_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	218 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_Update/ca
      -- CP-element group 225: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/type_cast_1412_Update/$exit
      -- 
    ca_3019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1412_inst_ack_1, ack => zeropad3D_CP_676_elements(225)); -- 
    -- CP-element group 226:  join  fork  transition  place  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	221 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	685 
    -- CP-element group 226: 	686 
    -- CP-element group 226: 	687 
    -- CP-element group 226: 	689 
    -- CP-element group 226:  members (16) 
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529
      -- CP-element group 226: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445__exit__
      -- CP-element group 226: 	 branch_block_stmt_223/assign_stmt_1400_to_assign_stmt_1445/$exit
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/$entry
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1448/$entry
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/$entry
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/$entry
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/$entry
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/$entry
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/SplitProtocol/$entry
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/SplitProtocol/Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/SplitProtocol/Sample/rr
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/SplitProtocol/Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/SplitProtocol/Update/cr
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1461/$entry
      -- CP-element group 226: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/$entry
      -- 
    rr_7463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(226), ack => type_cast_1458_inst_req_0); -- 
    cr_7468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(226), ack => type_cast_1458_inst_req_1); -- 
    zeropad3D_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(221) & zeropad3D_CP_676_elements(225);
      gj_zeropad3D_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	695 
    -- CP-element group 227: successors 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_Sample/ra
      -- CP-element group 227: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_sample_completed_
      -- 
    ra_3031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1472_inst_ack_0, ack => zeropad3D_CP_676_elements(227)); -- 
    -- CP-element group 228:  branch  transition  place  input  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	695 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (13) 
      -- CP-element group 228: 	 branch_block_stmt_223/if_stmt_1499__entry__
      -- CP-element group 228: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498__exit__
      -- CP-element group 228: 	 branch_block_stmt_223/R_orx_xcond1852_1500_place
      -- CP-element group 228: 	 branch_block_stmt_223/if_stmt_1499_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_223/if_stmt_1499_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_223/if_stmt_1499_else_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_223/if_stmt_1499_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_223/if_stmt_1499_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_223/if_stmt_1499_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_Update/ca
      -- CP-element group 228: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/$exit
      -- 
    ca_3036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1472_inst_ack_1, ack => zeropad3D_CP_676_elements(228)); -- 
    branch_req_3044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(228), ack => if_stmt_1499_branch_req_0); -- 
    -- CP-element group 229:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229: 	232 
    -- CP-element group 229:  members (18) 
      -- CP-element group 229: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535__entry__
      -- CP-element group 229: 	 branch_block_stmt_223/merge_stmt_1505__exit__
      -- CP-element group 229: 	 branch_block_stmt_223/whilex_xbody529_lorx_xlhsx_xfalse547
      -- CP-element group 229: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_Update/cr
      -- CP-element group 229: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/$entry
      -- CP-element group 229: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_223/if_stmt_1499_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_223/if_stmt_1499_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_Sample/rr
      -- CP-element group 229: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_update_start_
      -- CP-element group 229: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_223/merge_stmt_1505_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_223/whilex_xbody529_lorx_xlhsx_xfalse547_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_223/whilex_xbody529_lorx_xlhsx_xfalse547_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_223/merge_stmt_1505_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_223/merge_stmt_1505_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_223/merge_stmt_1505_PhiAck/dummy
      -- 
    if_choice_transition_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1499_branch_ack_1, ack => zeropad3D_CP_676_elements(229)); -- 
    cr_3071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(229), ack => type_cast_1509_inst_req_1); -- 
    rr_3066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(229), ack => type_cast_1509_inst_req_0); -- 
    -- CP-element group 230:  transition  place  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	696 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_223/whilex_xbody529_ifx_xthen565
      -- CP-element group 230: 	 branch_block_stmt_223/if_stmt_1499_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_223/if_stmt_1499_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_223/whilex_xbody529_ifx_xthen565_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_223/whilex_xbody529_ifx_xthen565_PhiReq/$exit
      -- 
    else_choice_transition_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1499_branch_ack_0, ack => zeropad3D_CP_676_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_Sample/ra
      -- CP-element group 231: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_sample_completed_
      -- 
    ra_3067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1509_inst_ack_0, ack => zeropad3D_CP_676_elements(231)); -- 
    -- CP-element group 232:  branch  transition  place  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	229 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (13) 
      -- CP-element group 232: 	 branch_block_stmt_223/if_stmt_1536_eval_test/$entry
      -- CP-element group 232: 	 branch_block_stmt_223/if_stmt_1536__entry__
      -- CP-element group 232: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535__exit__
      -- CP-element group 232: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_223/if_stmt_1536_eval_test/$exit
      -- CP-element group 232: 	 branch_block_stmt_223/if_stmt_1536_eval_test/branch_req
      -- CP-element group 232: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/$exit
      -- CP-element group 232: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_Update/ca
      -- CP-element group 232: 	 branch_block_stmt_223/if_stmt_1536_dead_link/$entry
      -- CP-element group 232: 	 branch_block_stmt_223/assign_stmt_1510_to_assign_stmt_1535/type_cast_1509_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_223/R_orx_xcond1853_1537_place
      -- CP-element group 232: 	 branch_block_stmt_223/if_stmt_1536_if_link/$entry
      -- CP-element group 232: 	 branch_block_stmt_223/if_stmt_1536_else_link/$entry
      -- 
    ca_3072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1509_inst_ack_1, ack => zeropad3D_CP_676_elements(232)); -- 
    branch_req_3080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(232), ack => if_stmt_1536_branch_req_0); -- 
    -- CP-element group 233:  fork  transition  place  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	249 
    -- CP-element group 233: 	250 
    -- CP-element group 233: 	252 
    -- CP-element group 233: 	254 
    -- CP-element group 233: 	256 
    -- CP-element group 233: 	258 
    -- CP-element group 233: 	260 
    -- CP-element group 233: 	262 
    -- CP-element group 233: 	264 
    -- CP-element group 233: 	267 
    -- CP-element group 233:  members (46) 
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705__entry__
      -- CP-element group 233: 	 branch_block_stmt_223/merge_stmt_1600__exit__
      -- CP-element group 233: 	 branch_block_stmt_223/if_stmt_1536_if_link/$exit
      -- CP-element group 233: 	 branch_block_stmt_223/if_stmt_1536_if_link/if_choice_transition
      -- CP-element group 233: 	 branch_block_stmt_223/lorx_xlhsx_xfalse547_ifx_xelse586
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_update_start_
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_Sample/rr
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_Update/cr
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_update_start_
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_Update/cr
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_update_start_
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_final_index_sum_regn_update_start
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_final_index_sum_regn_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_final_index_sum_regn_Update/req
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_complete/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_complete/req
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_update_start_
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/word_access_complete/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/word_access_complete/word_0/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/word_access_complete/word_0/cr
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_update_start_
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_Update/cr
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_update_start_
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_final_index_sum_regn_update_start
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_final_index_sum_regn_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_final_index_sum_regn_Update/req
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_complete/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_complete/req
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_update_start_
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Update/word_access_complete/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Update/word_access_complete/word_0/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Update/word_access_complete/word_0/cr
      -- CP-element group 233: 	 branch_block_stmt_223/merge_stmt_1600_PhiReqMerge
      -- CP-element group 233: 	 branch_block_stmt_223/lorx_xlhsx_xfalse547_ifx_xelse586_PhiReq/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/lorx_xlhsx_xfalse547_ifx_xelse586_PhiReq/$exit
      -- CP-element group 233: 	 branch_block_stmt_223/merge_stmt_1600_PhiAck/$entry
      -- CP-element group 233: 	 branch_block_stmt_223/merge_stmt_1600_PhiAck/$exit
      -- CP-element group 233: 	 branch_block_stmt_223/merge_stmt_1600_PhiAck/dummy
      -- 
    if_choice_transition_3085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1536_branch_ack_1, ack => zeropad3D_CP_676_elements(233)); -- 
    rr_3243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => type_cast_1604_inst_req_0); -- 
    cr_3248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => type_cast_1604_inst_req_1); -- 
    cr_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => type_cast_1668_inst_req_1); -- 
    req_3293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => array_obj_ref_1674_index_offset_req_1); -- 
    req_3308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => addr_of_1675_final_reg_req_1); -- 
    cr_3353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => ptr_deref_1679_load_0_req_1); -- 
    cr_3372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => type_cast_1693_inst_req_1); -- 
    req_3403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => array_obj_ref_1699_index_offset_req_1); -- 
    req_3418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => addr_of_1700_final_reg_req_1); -- 
    cr_3468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(233), ack => ptr_deref_1703_store_0_req_1); -- 
    -- CP-element group 234:  transition  place  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	696 
    -- CP-element group 234:  members (5) 
      -- CP-element group 234: 	 branch_block_stmt_223/if_stmt_1536_else_link/$exit
      -- CP-element group 234: 	 branch_block_stmt_223/if_stmt_1536_else_link/else_choice_transition
      -- CP-element group 234: 	 branch_block_stmt_223/lorx_xlhsx_xfalse547_ifx_xthen565
      -- CP-element group 234: 	 branch_block_stmt_223/lorx_xlhsx_xfalse547_ifx_xthen565_PhiReq/$entry
      -- CP-element group 234: 	 branch_block_stmt_223/lorx_xlhsx_xfalse547_ifx_xthen565_PhiReq/$exit
      -- 
    else_choice_transition_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1536_branch_ack_0, ack => zeropad3D_CP_676_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	696 
    -- CP-element group 235: successors 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_Sample/ra
      -- 
    ra_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1546_inst_ack_0, ack => zeropad3D_CP_676_elements(235)); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	696 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	239 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_Update/ca
      -- 
    ca_3108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1546_inst_ack_1, ack => zeropad3D_CP_676_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	696 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_Sample/ra
      -- 
    ra_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1551_inst_ack_0, ack => zeropad3D_CP_676_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	696 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_Update/ca
      -- 
    ca_3122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1551_inst_ack_1, ack => zeropad3D_CP_676_elements(238)); -- 
    -- CP-element group 239:  join  transition  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	236 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_Sample/rr
      -- 
    rr_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(239), ack => type_cast_1585_inst_req_0); -- 
    zeropad3D_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(236) & zeropad3D_CP_676_elements(238);
      gj_zeropad3D_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_sample_completed_
      -- CP-element group 240: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_Sample/ra
      -- 
    ra_3131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1585_inst_ack_0, ack => zeropad3D_CP_676_elements(240)); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	696 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (16) 
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_update_completed_
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_Update/ca
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_resized_1
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_scaled_1
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_computed_1
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_resize_1/$entry
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_resize_1/$exit
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_resize_1/index_resize_req
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_resize_1/index_resize_ack
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_scale_1/$entry
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_scale_1/$exit
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_scale_1/scale_rename_req
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_index_scale_1/scale_rename_ack
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_final_index_sum_regn_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_final_index_sum_regn_Sample/req
      -- 
    ca_3136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1585_inst_ack_1, ack => zeropad3D_CP_676_elements(241)); -- 
    req_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(241), ack => array_obj_ref_1591_index_offset_req_0); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	248 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_final_index_sum_regn_sample_complete
      -- CP-element group 242: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_final_index_sum_regn_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_final_index_sum_regn_Sample/ack
      -- 
    ack_3162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1591_index_offset_ack_0, ack => zeropad3D_CP_676_elements(242)); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	696 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (11) 
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_root_address_calculated
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_offset_calculated
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_final_index_sum_regn_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_final_index_sum_regn_Update/ack
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_base_plus_offset/$entry
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_base_plus_offset/$exit
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_base_plus_offset/sum_rename_req
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_base_plus_offset/sum_rename_ack
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_request/$entry
      -- CP-element group 243: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_request/req
      -- 
    ack_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1591_index_offset_ack_1, ack => zeropad3D_CP_676_elements(243)); -- 
    req_3176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(243), ack => addr_of_1592_final_reg_req_0); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_request/$exit
      -- CP-element group 244: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_request/ack
      -- 
    ack_3177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1592_final_reg_ack_0, ack => zeropad3D_CP_676_elements(244)); -- 
    -- CP-element group 245:  join  fork  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	696 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (28) 
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_complete/$exit
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_complete/ack
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_base_address_calculated
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_word_address_calculated
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_root_address_calculated
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_base_address_resized
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_base_addr_resize/$entry
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_base_addr_resize/$exit
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_base_addr_resize/base_resize_req
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_base_addr_resize/base_resize_ack
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_base_plus_offset/$entry
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_base_plus_offset/$exit
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_base_plus_offset/sum_rename_req
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_base_plus_offset/sum_rename_ack
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_word_addrgen/$entry
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_word_addrgen/$exit
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_word_addrgen/root_register_req
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_word_addrgen/root_register_ack
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/ptr_deref_1595_Split/$entry
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/ptr_deref_1595_Split/$exit
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/ptr_deref_1595_Split/split_req
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/ptr_deref_1595_Split/split_ack
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/word_access_start/$entry
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/word_access_start/word_0/$entry
      -- CP-element group 245: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/word_access_start/word_0/rr
      -- 
    ack_3182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1592_final_reg_ack_1, ack => zeropad3D_CP_676_elements(245)); -- 
    rr_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(245), ack => ptr_deref_1595_store_0_req_0); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (5) 
      -- CP-element group 246: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/word_access_start/$exit
      -- CP-element group 246: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/word_access_start/word_0/$exit
      -- CP-element group 246: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Sample/word_access_start/word_0/ra
      -- 
    ra_3221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1595_store_0_ack_0, ack => zeropad3D_CP_676_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	696 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (5) 
      -- CP-element group 247: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Update/word_access_complete/$exit
      -- CP-element group 247: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Update/word_access_complete/word_0/$exit
      -- CP-element group 247: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Update/word_access_complete/word_0/ca
      -- 
    ca_3232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1595_store_0_ack_1, ack => zeropad3D_CP_676_elements(247)); -- 
    -- CP-element group 248:  join  transition  place  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	242 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	697 
    -- CP-element group 248:  members (5) 
      -- CP-element group 248: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598__exit__
      -- CP-element group 248: 	 branch_block_stmt_223/ifx_xthen565_ifx_xend634
      -- CP-element group 248: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/$exit
      -- CP-element group 248: 	 branch_block_stmt_223/ifx_xthen565_ifx_xend634_PhiReq/$entry
      -- CP-element group 248: 	 branch_block_stmt_223/ifx_xthen565_ifx_xend634_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(242) & zeropad3D_CP_676_elements(247);
      gj_zeropad3D_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	233 
    -- CP-element group 249: successors 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_Sample/ra
      -- 
    ra_3244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1604_inst_ack_0, ack => zeropad3D_CP_676_elements(249)); -- 
    -- CP-element group 250:  fork  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	233 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250: 	259 
    -- CP-element group 250:  members (9) 
      -- CP-element group 250: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1604_Update/ca
      -- CP-element group 250: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_Sample/rr
      -- CP-element group 250: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_Sample/rr
      -- 
    ca_3249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1604_inst_ack_1, ack => zeropad3D_CP_676_elements(250)); -- 
    rr_3257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(250), ack => type_cast_1668_inst_req_0); -- 
    rr_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(250), ack => type_cast_1693_inst_req_0); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_Sample/ra
      -- 
    ra_3258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1668_inst_ack_0, ack => zeropad3D_CP_676_elements(251)); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	233 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (16) 
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1668_Update/ca
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_resized_1
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_scaled_1
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_computed_1
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_resize_1/$entry
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_resize_1/$exit
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_resize_1/index_resize_req
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_resize_1/index_resize_ack
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_scale_1/$entry
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_scale_1/$exit
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_scale_1/scale_rename_req
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_index_scale_1/scale_rename_ack
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_final_index_sum_regn_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_final_index_sum_regn_Sample/req
      -- 
    ca_3263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1668_inst_ack_1, ack => zeropad3D_CP_676_elements(252)); -- 
    req_3288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(252), ack => array_obj_ref_1674_index_offset_req_0); -- 
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	268 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_final_index_sum_regn_sample_complete
      -- CP-element group 253: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_final_index_sum_regn_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_final_index_sum_regn_Sample/ack
      -- 
    ack_3289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1674_index_offset_ack_0, ack => zeropad3D_CP_676_elements(253)); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	233 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (11) 
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_root_address_calculated
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_offset_calculated
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_final_index_sum_regn_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_final_index_sum_regn_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_base_plus_offset/$entry
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_base_plus_offset/$exit
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_base_plus_offset/sum_rename_req
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1674_base_plus_offset/sum_rename_ack
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_request/$entry
      -- CP-element group 254: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_request/req
      -- 
    ack_3294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1674_index_offset_ack_1, ack => zeropad3D_CP_676_elements(254)); -- 
    req_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(254), ack => addr_of_1675_final_reg_req_0); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_request/$exit
      -- CP-element group 255: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_request/ack
      -- 
    ack_3304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1675_final_reg_ack_0, ack => zeropad3D_CP_676_elements(255)); -- 
    -- CP-element group 256:  join  fork  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	233 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (24) 
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_complete/$exit
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1675_complete/ack
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_base_address_calculated
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_word_address_calculated
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_root_address_calculated
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_base_address_resized
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_base_addr_resize/$entry
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_base_addr_resize/$exit
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_base_addr_resize/base_resize_req
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_base_addr_resize/base_resize_ack
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_base_plus_offset/$entry
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_base_plus_offset/$exit
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_base_plus_offset/sum_rename_req
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_base_plus_offset/sum_rename_ack
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_word_addrgen/$entry
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_word_addrgen/$exit
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_word_addrgen/root_register_req
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_word_addrgen/root_register_ack
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Sample/word_access_start/$entry
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Sample/word_access_start/word_0/$entry
      -- CP-element group 256: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Sample/word_access_start/word_0/rr
      -- 
    ack_3309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1675_final_reg_ack_1, ack => zeropad3D_CP_676_elements(256)); -- 
    rr_3342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(256), ack => ptr_deref_1679_load_0_req_0); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257:  members (5) 
      -- CP-element group 257: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Sample/word_access_start/$exit
      -- CP-element group 257: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Sample/word_access_start/word_0/$exit
      -- CP-element group 257: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Sample/word_access_start/word_0/ra
      -- 
    ra_3343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1679_load_0_ack_0, ack => zeropad3D_CP_676_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	233 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	265 
    -- CP-element group 258:  members (9) 
      -- CP-element group 258: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/word_access_complete/$exit
      -- CP-element group 258: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/word_access_complete/word_0/$exit
      -- CP-element group 258: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/word_access_complete/word_0/ca
      -- CP-element group 258: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/ptr_deref_1679_Merge/$entry
      -- CP-element group 258: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/ptr_deref_1679_Merge/$exit
      -- CP-element group 258: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/ptr_deref_1679_Merge/merge_req
      -- CP-element group 258: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1679_Update/ptr_deref_1679_Merge/merge_ack
      -- 
    ca_3354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1679_load_0_ack_1, ack => zeropad3D_CP_676_elements(258)); -- 
    -- CP-element group 259:  transition  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	250 
    -- CP-element group 259: successors 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_sample_completed_
      -- CP-element group 259: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_Sample/ra
      -- 
    ra_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1693_inst_ack_0, ack => zeropad3D_CP_676_elements(259)); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	233 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (16) 
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/type_cast_1693_Update/ca
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_resized_1
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_scaled_1
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_computed_1
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_resize_1/$entry
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_resize_1/$exit
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_resize_1/index_resize_req
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_resize_1/index_resize_ack
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_scale_1/$entry
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_scale_1/$exit
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_scale_1/scale_rename_req
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_index_scale_1/scale_rename_ack
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_final_index_sum_regn_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_final_index_sum_regn_Sample/req
      -- 
    ca_3373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1693_inst_ack_1, ack => zeropad3D_CP_676_elements(260)); -- 
    req_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(260), ack => array_obj_ref_1699_index_offset_req_0); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	268 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_final_index_sum_regn_sample_complete
      -- CP-element group 261: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_final_index_sum_regn_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_final_index_sum_regn_Sample/ack
      -- 
    ack_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1699_index_offset_ack_0, ack => zeropad3D_CP_676_elements(261)); -- 
    -- CP-element group 262:  transition  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	233 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (11) 
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_root_address_calculated
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_offset_calculated
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_final_index_sum_regn_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_final_index_sum_regn_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_base_plus_offset/$entry
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_base_plus_offset/$exit
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_base_plus_offset/sum_rename_req
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/array_obj_ref_1699_base_plus_offset/sum_rename_ack
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_request/$entry
      -- CP-element group 262: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_request/req
      -- 
    ack_3404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1699_index_offset_ack_1, ack => zeropad3D_CP_676_elements(262)); -- 
    req_3413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(262), ack => addr_of_1700_final_reg_req_0); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_request/$exit
      -- CP-element group 263: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_request/ack
      -- 
    ack_3414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1700_final_reg_ack_0, ack => zeropad3D_CP_676_elements(263)); -- 
    -- CP-element group 264:  fork  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	233 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (19) 
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_complete/$exit
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/addr_of_1700_complete/ack
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_base_address_calculated
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_word_address_calculated
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_root_address_calculated
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_base_address_resized
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_base_addr_resize/$entry
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_base_addr_resize/$exit
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_base_addr_resize/base_resize_req
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_base_addr_resize/base_resize_ack
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_base_plus_offset/$entry
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_base_plus_offset/$exit
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_base_plus_offset/sum_rename_req
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_base_plus_offset/sum_rename_ack
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_word_addrgen/$entry
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_word_addrgen/$exit
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_word_addrgen/root_register_req
      -- CP-element group 264: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_word_addrgen/root_register_ack
      -- 
    ack_3419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1700_final_reg_ack_1, ack => zeropad3D_CP_676_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	258 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (9) 
      -- CP-element group 265: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/ptr_deref_1703_Split/$entry
      -- CP-element group 265: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/ptr_deref_1703_Split/$exit
      -- CP-element group 265: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/ptr_deref_1703_Split/split_req
      -- CP-element group 265: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/ptr_deref_1703_Split/split_ack
      -- CP-element group 265: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/word_access_start/$entry
      -- CP-element group 265: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/word_access_start/word_0/$entry
      -- CP-element group 265: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/word_access_start/word_0/rr
      -- 
    rr_3457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(265), ack => ptr_deref_1703_store_0_req_0); -- 
    zeropad3D_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(258) & zeropad3D_CP_676_elements(264);
      gj_zeropad3D_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266:  members (5) 
      -- CP-element group 266: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/word_access_start/$exit
      -- CP-element group 266: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/word_access_start/word_0/$exit
      -- CP-element group 266: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Sample/word_access_start/word_0/ra
      -- 
    ra_3458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1703_store_0_ack_0, ack => zeropad3D_CP_676_elements(266)); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	233 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (5) 
      -- CP-element group 267: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Update/word_access_complete/$exit
      -- CP-element group 267: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Update/word_access_complete/word_0/$exit
      -- CP-element group 267: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/ptr_deref_1703_Update/word_access_complete/word_0/ca
      -- 
    ca_3469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1703_store_0_ack_1, ack => zeropad3D_CP_676_elements(267)); -- 
    -- CP-element group 268:  join  transition  place  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	253 
    -- CP-element group 268: 	261 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	697 
    -- CP-element group 268:  members (5) 
      -- CP-element group 268: 	 branch_block_stmt_223/ifx_xelse586_ifx_xend634
      -- CP-element group 268: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705__exit__
      -- CP-element group 268: 	 branch_block_stmt_223/assign_stmt_1605_to_assign_stmt_1705/$exit
      -- CP-element group 268: 	 branch_block_stmt_223/ifx_xelse586_ifx_xend634_PhiReq/$entry
      -- CP-element group 268: 	 branch_block_stmt_223/ifx_xelse586_ifx_xend634_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(253) & zeropad3D_CP_676_elements(261) & zeropad3D_CP_676_elements(267);
      gj_zeropad3D_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	697 
    -- CP-element group 269: successors 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_sample_completed_
      -- CP-element group 269: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_Sample/ra
      -- 
    ra_3481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1711_inst_ack_0, ack => zeropad3D_CP_676_elements(269)); -- 
    -- CP-element group 270:  branch  transition  place  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	697 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (13) 
      -- CP-element group 270: 	 branch_block_stmt_223/if_stmt_1726__entry__
      -- CP-element group 270: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725__exit__
      -- CP-element group 270: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/$exit
      -- CP-element group 270: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_update_completed_
      -- CP-element group 270: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_Update/ca
      -- CP-element group 270: 	 branch_block_stmt_223/if_stmt_1726_dead_link/$entry
      -- CP-element group 270: 	 branch_block_stmt_223/if_stmt_1726_eval_test/$entry
      -- CP-element group 270: 	 branch_block_stmt_223/if_stmt_1726_eval_test/$exit
      -- CP-element group 270: 	 branch_block_stmt_223/if_stmt_1726_eval_test/branch_req
      -- CP-element group 270: 	 branch_block_stmt_223/R_cmp642_1727_place
      -- CP-element group 270: 	 branch_block_stmt_223/if_stmt_1726_if_link/$entry
      -- CP-element group 270: 	 branch_block_stmt_223/if_stmt_1726_else_link/$entry
      -- 
    ca_3486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1711_inst_ack_1, ack => zeropad3D_CP_676_elements(270)); -- 
    branch_req_3494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(270), ack => if_stmt_1726_branch_req_0); -- 
    -- CP-element group 271:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	706 
    -- CP-element group 271: 	707 
    -- CP-element group 271: 	709 
    -- CP-element group 271: 	710 
    -- CP-element group 271: 	712 
    -- CP-element group 271: 	713 
    -- CP-element group 271:  members (40) 
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686
      -- CP-element group 271: 	 branch_block_stmt_223/assign_stmt_1738__exit__
      -- CP-element group 271: 	 branch_block_stmt_223/assign_stmt_1738__entry__
      -- CP-element group 271: 	 branch_block_stmt_223/merge_stmt_1732__exit__
      -- CP-element group 271: 	 branch_block_stmt_223/if_stmt_1726_if_link/$exit
      -- CP-element group 271: 	 branch_block_stmt_223/if_stmt_1726_if_link/if_choice_transition
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xend634_ifx_xthen644
      -- CP-element group 271: 	 branch_block_stmt_223/assign_stmt_1738/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/assign_stmt_1738/$exit
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xend634_ifx_xthen644_PhiReq/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xend634_ifx_xthen644_PhiReq/$exit
      -- CP-element group 271: 	 branch_block_stmt_223/merge_stmt_1732_PhiReqMerge
      -- CP-element group 271: 	 branch_block_stmt_223/merge_stmt_1732_PhiAck/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/merge_stmt_1732_PhiAck/$exit
      -- CP-element group 271: 	 branch_block_stmt_223/merge_stmt_1732_PhiAck/dummy
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/SplitProtocol/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/SplitProtocol/Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/SplitProtocol/Sample/rr
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/SplitProtocol/Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/SplitProtocol/Update/cr
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Sample/rr
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Update/cr
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Sample/rr
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1726_branch_ack_1, ack => zeropad3D_CP_676_elements(271)); -- 
    rr_7631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(271), ack => type_cast_1806_inst_req_0); -- 
    cr_7636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(271), ack => type_cast_1806_inst_req_1); -- 
    rr_7654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(271), ack => type_cast_1800_inst_req_0); -- 
    cr_7659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(271), ack => type_cast_1800_inst_req_1); -- 
    rr_7677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(271), ack => type_cast_1793_inst_req_0); -- 
    cr_7682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(271), ack => type_cast_1793_inst_req_1); -- 
    -- CP-element group 272:  fork  transition  place  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272: 	274 
    -- CP-element group 272: 	276 
    -- CP-element group 272: 	278 
    -- CP-element group 272:  members (24) 
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782__entry__
      -- CP-element group 272: 	 branch_block_stmt_223/merge_stmt_1740__exit__
      -- CP-element group 272: 	 branch_block_stmt_223/if_stmt_1726_else_link/$exit
      -- CP-element group 272: 	 branch_block_stmt_223/if_stmt_1726_else_link/else_choice_transition
      -- CP-element group 272: 	 branch_block_stmt_223/ifx_xend634_ifx_xelse649
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/$entry
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_update_start_
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_update_start_
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_update_start_
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_223/ifx_xend634_ifx_xelse649_PhiReq/$entry
      -- CP-element group 272: 	 branch_block_stmt_223/ifx_xend634_ifx_xelse649_PhiReq/$exit
      -- CP-element group 272: 	 branch_block_stmt_223/merge_stmt_1740_PhiReqMerge
      -- CP-element group 272: 	 branch_block_stmt_223/merge_stmt_1740_PhiAck/$entry
      -- CP-element group 272: 	 branch_block_stmt_223/merge_stmt_1740_PhiAck/$exit
      -- CP-element group 272: 	 branch_block_stmt_223/merge_stmt_1740_PhiAck/dummy
      -- 
    else_choice_transition_3503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1726_branch_ack_0, ack => zeropad3D_CP_676_elements(272)); -- 
    rr_3519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(272), ack => type_cast_1750_inst_req_0); -- 
    cr_3524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(272), ack => type_cast_1750_inst_req_1); -- 
    cr_3538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(272), ack => type_cast_1759_inst_req_1); -- 
    cr_3552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(272), ack => type_cast_1776_inst_req_1); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_Sample/ra
      -- 
    ra_3520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1750_inst_ack_0, ack => zeropad3D_CP_676_elements(273)); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1750_Update/ca
      -- CP-element group 274: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_Sample/rr
      -- 
    ca_3525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1750_inst_ack_1, ack => zeropad3D_CP_676_elements(274)); -- 
    rr_3533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(274), ack => type_cast_1759_inst_req_0); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_sample_completed_
      -- CP-element group 275: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_Sample/ra
      -- 
    ra_3534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1759_inst_ack_0, ack => zeropad3D_CP_676_elements(275)); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	272 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1759_Update/ca
      -- CP-element group 276: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_Sample/rr
      -- 
    ca_3539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1759_inst_ack_1, ack => zeropad3D_CP_676_elements(276)); -- 
    rr_3547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(276), ack => type_cast_1776_inst_req_0); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_sample_completed_
      -- CP-element group 277: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_Sample/ra
      -- 
    ra_3548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1776_inst_ack_0, ack => zeropad3D_CP_676_elements(277)); -- 
    -- CP-element group 278:  branch  transition  place  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	272 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (13) 
      -- CP-element group 278: 	 branch_block_stmt_223/if_stmt_1783__entry__
      -- CP-element group 278: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782__exit__
      -- CP-element group 278: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/$exit
      -- CP-element group 278: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_223/assign_stmt_1746_to_assign_stmt_1782/type_cast_1776_Update/ca
      -- CP-element group 278: 	 branch_block_stmt_223/if_stmt_1783_dead_link/$entry
      -- CP-element group 278: 	 branch_block_stmt_223/if_stmt_1783_eval_test/$entry
      -- CP-element group 278: 	 branch_block_stmt_223/if_stmt_1783_eval_test/$exit
      -- CP-element group 278: 	 branch_block_stmt_223/if_stmt_1783_eval_test/branch_req
      -- CP-element group 278: 	 branch_block_stmt_223/R_cmp677_1784_place
      -- CP-element group 278: 	 branch_block_stmt_223/if_stmt_1783_if_link/$entry
      -- CP-element group 278: 	 branch_block_stmt_223/if_stmt_1783_else_link/$entry
      -- 
    ca_3553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1776_inst_ack_1, ack => zeropad3D_CP_676_elements(278)); -- 
    branch_req_3561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(278), ack => if_stmt_1783_branch_req_0); -- 
    -- CP-element group 279:  fork  transition  place  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279: 	282 
    -- CP-element group 279: 	284 
    -- CP-element group 279:  members (27) 
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844__entry__
      -- CP-element group 279: 	 branch_block_stmt_223/merge_stmt_1811__exit__
      -- CP-element group 279: 	 branch_block_stmt_223/if_stmt_1783_if_link/$exit
      -- CP-element group 279: 	 branch_block_stmt_223/if_stmt_1783_if_link/if_choice_transition
      -- CP-element group 279: 	 branch_block_stmt_223/ifx_xelse649_whilex_xend687
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/$entry
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_sample_start_
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_update_start_
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_word_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_root_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Sample/word_access_start/$entry
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Sample/word_access_start/word_0/$entry
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Sample/word_access_start/word_0/rr
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/word_access_complete/$entry
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/word_access_complete/word_0/$entry
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/word_access_complete/word_0/cr
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_update_start_
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_Update/cr
      -- CP-element group 279: 	 branch_block_stmt_223/ifx_xelse649_whilex_xend687_PhiReq/$entry
      -- CP-element group 279: 	 branch_block_stmt_223/ifx_xelse649_whilex_xend687_PhiReq/$exit
      -- CP-element group 279: 	 branch_block_stmt_223/merge_stmt_1811_PhiReqMerge
      -- CP-element group 279: 	 branch_block_stmt_223/merge_stmt_1811_PhiAck/$entry
      -- CP-element group 279: 	 branch_block_stmt_223/merge_stmt_1811_PhiAck/$exit
      -- CP-element group 279: 	 branch_block_stmt_223/merge_stmt_1811_PhiAck/dummy
      -- 
    if_choice_transition_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1783_branch_ack_1, ack => zeropad3D_CP_676_elements(279)); -- 
    rr_3591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(279), ack => LOAD_pad_1813_load_0_req_0); -- 
    cr_3602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(279), ack => LOAD_pad_1813_load_0_req_1); -- 
    cr_3621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(279), ack => type_cast_1817_inst_req_1); -- 
    -- CP-element group 280:  fork  transition  place  input  output  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	698 
    -- CP-element group 280: 	699 
    -- CP-element group 280: 	701 
    -- CP-element group 280: 	702 
    -- CP-element group 280: 	704 
    -- CP-element group 280:  members (22) 
      -- CP-element group 280: 	 branch_block_stmt_223/if_stmt_1783_else_link/$exit
      -- CP-element group 280: 	 branch_block_stmt_223/if_stmt_1783_else_link/else_choice_transition
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/SplitProtocol/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/SplitProtocol/Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/SplitProtocol/Sample/rr
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/SplitProtocol/Update/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/SplitProtocol/Update/cr
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Sample/rr
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Update/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Update/cr
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1790/$entry
      -- CP-element group 280: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/$entry
      -- 
    else_choice_transition_3570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1783_branch_ack_0, ack => zeropad3D_CP_676_elements(280)); -- 
    rr_7574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(280), ack => type_cast_1808_inst_req_0); -- 
    cr_7579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(280), ack => type_cast_1808_inst_req_1); -- 
    rr_7597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(280), ack => type_cast_1802_inst_req_0); -- 
    cr_7602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(280), ack => type_cast_1802_inst_req_1); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (5) 
      -- CP-element group 281: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Sample/word_access_start/$exit
      -- CP-element group 281: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Sample/word_access_start/word_0/$exit
      -- CP-element group 281: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Sample/word_access_start/word_0/ra
      -- 
    ra_3592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1813_load_0_ack_0, ack => zeropad3D_CP_676_elements(281)); -- 
    -- CP-element group 282:  transition  input  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	279 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (12) 
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/word_access_complete/$exit
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/word_access_complete/word_0/$exit
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/word_access_complete/word_0/ca
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/LOAD_pad_1813_Merge/$entry
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/LOAD_pad_1813_Merge/$exit
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/LOAD_pad_1813_Merge/merge_req
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/LOAD_pad_1813_Update/LOAD_pad_1813_Merge/merge_ack
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_sample_start_
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_Sample/rr
      -- 
    ca_3603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_1813_load_0_ack_1, ack => zeropad3D_CP_676_elements(282)); -- 
    rr_3616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(282), ack => type_cast_1817_inst_req_0); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_sample_completed_
      -- CP-element group 283: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_Sample/ra
      -- 
    ra_3617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1817_inst_ack_0, ack => zeropad3D_CP_676_elements(283)); -- 
    -- CP-element group 284:  fork  transition  place  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	279 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	731 
    -- CP-element group 284: 	732 
    -- CP-element group 284: 	734 
    -- CP-element group 284: 	735 
    -- CP-element group 284: 	737 
    -- CP-element group 284:  members (25) 
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751
      -- CP-element group 284: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844__exit__
      -- CP-element group 284: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/$exit
      -- CP-element group 284: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_update_completed_
      -- CP-element group 284: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_223/assign_stmt_1814_to_assign_stmt_1844/type_cast_1817_Update/ca
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/SplitProtocol/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/SplitProtocol/Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/SplitProtocol/Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/SplitProtocol/Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/SplitProtocol/Update/cr
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/SplitProtocol/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/SplitProtocol/Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/SplitProtocol/Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/SplitProtocol/Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/SplitProtocol/Update/cr
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1847/$entry
      -- CP-element group 284: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/$entry
      -- 
    ca_3622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1817_inst_ack_1, ack => zeropad3D_CP_676_elements(284)); -- 
    rr_7790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(284), ack => type_cast_1865_inst_req_0); -- 
    cr_7795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(284), ack => type_cast_1865_inst_req_1); -- 
    rr_7813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(284), ack => type_cast_1859_inst_req_0); -- 
    cr_7818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(284), ack => type_cast_1859_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	743 
    -- CP-element group 285: successors 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_Sample/ra
      -- 
    ra_3634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1870_inst_ack_0, ack => zeropad3D_CP_676_elements(285)); -- 
    -- CP-element group 286:  branch  transition  place  input  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	743 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (13) 
      -- CP-element group 286: 	 branch_block_stmt_223/if_stmt_1897__entry__
      -- CP-element group 286: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896__exit__
      -- CP-element group 286: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/$exit
      -- CP-element group 286: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_Update/ca
      -- CP-element group 286: 	 branch_block_stmt_223/if_stmt_1897_dead_link/$entry
      -- CP-element group 286: 	 branch_block_stmt_223/if_stmt_1897_eval_test/$entry
      -- CP-element group 286: 	 branch_block_stmt_223/if_stmt_1897_eval_test/$exit
      -- CP-element group 286: 	 branch_block_stmt_223/if_stmt_1897_eval_test/branch_req
      -- CP-element group 286: 	 branch_block_stmt_223/R_orx_xcond1854_1898_place
      -- CP-element group 286: 	 branch_block_stmt_223/if_stmt_1897_if_link/$entry
      -- CP-element group 286: 	 branch_block_stmt_223/if_stmt_1897_else_link/$entry
      -- 
    ca_3639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1870_inst_ack_1, ack => zeropad3D_CP_676_elements(286)); -- 
    branch_req_3647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(286), ack => if_stmt_1897_branch_req_0); -- 
    -- CP-element group 287:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	289 
    -- CP-element group 287: 	290 
    -- CP-element group 287:  members (18) 
      -- CP-element group 287: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933__entry__
      -- CP-element group 287: 	 branch_block_stmt_223/merge_stmt_1903__exit__
      -- CP-element group 287: 	 branch_block_stmt_223/if_stmt_1897_if_link/$exit
      -- CP-element group 287: 	 branch_block_stmt_223/if_stmt_1897_if_link/if_choice_transition
      -- CP-element group 287: 	 branch_block_stmt_223/whilex_xbody751_lorx_xlhsx_xfalse769
      -- CP-element group 287: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/$entry
      -- CP-element group 287: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_update_start_
      -- CP-element group 287: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_Sample/rr
      -- CP-element group 287: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_Update/cr
      -- CP-element group 287: 	 branch_block_stmt_223/whilex_xbody751_lorx_xlhsx_xfalse769_PhiReq/$entry
      -- CP-element group 287: 	 branch_block_stmt_223/whilex_xbody751_lorx_xlhsx_xfalse769_PhiReq/$exit
      -- CP-element group 287: 	 branch_block_stmt_223/merge_stmt_1903_PhiReqMerge
      -- CP-element group 287: 	 branch_block_stmt_223/merge_stmt_1903_PhiAck/$entry
      -- CP-element group 287: 	 branch_block_stmt_223/merge_stmt_1903_PhiAck/$exit
      -- CP-element group 287: 	 branch_block_stmt_223/merge_stmt_1903_PhiAck/dummy
      -- 
    if_choice_transition_3652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1897_branch_ack_1, ack => zeropad3D_CP_676_elements(287)); -- 
    rr_3669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(287), ack => type_cast_1907_inst_req_0); -- 
    cr_3674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(287), ack => type_cast_1907_inst_req_1); -- 
    -- CP-element group 288:  transition  place  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	744 
    -- CP-element group 288:  members (5) 
      -- CP-element group 288: 	 branch_block_stmt_223/if_stmt_1897_else_link/$exit
      -- CP-element group 288: 	 branch_block_stmt_223/if_stmt_1897_else_link/else_choice_transition
      -- CP-element group 288: 	 branch_block_stmt_223/whilex_xbody751_ifx_xthen786
      -- CP-element group 288: 	 branch_block_stmt_223/whilex_xbody751_ifx_xthen786_PhiReq/$entry
      -- CP-element group 288: 	 branch_block_stmt_223/whilex_xbody751_ifx_xthen786_PhiReq/$exit
      -- 
    else_choice_transition_3656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1897_branch_ack_0, ack => zeropad3D_CP_676_elements(288)); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	287 
    -- CP-element group 289: successors 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_sample_completed_
      -- CP-element group 289: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_Sample/ra
      -- 
    ra_3670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1907_inst_ack_0, ack => zeropad3D_CP_676_elements(289)); -- 
    -- CP-element group 290:  branch  transition  place  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	287 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (13) 
      -- CP-element group 290: 	 branch_block_stmt_223/if_stmt_1934__entry__
      -- CP-element group 290: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933__exit__
      -- CP-element group 290: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/$exit
      -- CP-element group 290: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_223/assign_stmt_1908_to_assign_stmt_1933/type_cast_1907_Update/ca
      -- CP-element group 290: 	 branch_block_stmt_223/if_stmt_1934_dead_link/$entry
      -- CP-element group 290: 	 branch_block_stmt_223/if_stmt_1934_eval_test/$entry
      -- CP-element group 290: 	 branch_block_stmt_223/if_stmt_1934_eval_test/$exit
      -- CP-element group 290: 	 branch_block_stmt_223/if_stmt_1934_eval_test/branch_req
      -- CP-element group 290: 	 branch_block_stmt_223/R_orx_xcond1855_1935_place
      -- CP-element group 290: 	 branch_block_stmt_223/if_stmt_1934_if_link/$entry
      -- CP-element group 290: 	 branch_block_stmt_223/if_stmt_1934_else_link/$entry
      -- 
    ca_3675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1907_inst_ack_1, ack => zeropad3D_CP_676_elements(290)); -- 
    branch_req_3683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(290), ack => if_stmt_1934_branch_req_0); -- 
    -- CP-element group 291:  fork  transition  place  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	307 
    -- CP-element group 291: 	308 
    -- CP-element group 291: 	310 
    -- CP-element group 291: 	312 
    -- CP-element group 291: 	314 
    -- CP-element group 291: 	316 
    -- CP-element group 291: 	318 
    -- CP-element group 291: 	320 
    -- CP-element group 291: 	322 
    -- CP-element group 291: 	325 
    -- CP-element group 291:  members (46) 
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103__entry__
      -- CP-element group 291: 	 branch_block_stmt_223/merge_stmt_1998__exit__
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_Update/cr
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/word_access_complete/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_complete/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/word_access_complete/word_0/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_update_start_
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_update_start_
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/word_access_complete/word_0/cr
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_final_index_sum_regn_Update/req
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_final_index_sum_regn_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Update/word_access_complete/word_0/cr
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_final_index_sum_regn_update_start
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Update/word_access_complete/word_0/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_update_start_
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Update/word_access_complete/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_update_start_
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_complete/req
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_complete/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_Update/cr
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_update_start_
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_update_start_
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_Sample/rr
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_final_index_sum_regn_Update/req
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_final_index_sum_regn_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_final_index_sum_regn_update_start
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_Update/cr
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_Sample/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_update_start_
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_complete/req
      -- CP-element group 291: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_sample_start_
      -- CP-element group 291: 	 branch_block_stmt_223/if_stmt_1934_if_link/$exit
      -- CP-element group 291: 	 branch_block_stmt_223/if_stmt_1934_if_link/if_choice_transition
      -- CP-element group 291: 	 branch_block_stmt_223/lorx_xlhsx_xfalse769_ifx_xelse807
      -- CP-element group 291: 	 branch_block_stmt_223/lorx_xlhsx_xfalse769_ifx_xelse807_PhiReq/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/lorx_xlhsx_xfalse769_ifx_xelse807_PhiReq/$exit
      -- CP-element group 291: 	 branch_block_stmt_223/merge_stmt_1998_PhiReqMerge
      -- CP-element group 291: 	 branch_block_stmt_223/merge_stmt_1998_PhiAck/$entry
      -- CP-element group 291: 	 branch_block_stmt_223/merge_stmt_1998_PhiAck/$exit
      -- CP-element group 291: 	 branch_block_stmt_223/merge_stmt_1998_PhiAck/dummy
      -- 
    if_choice_transition_3688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1934_branch_ack_1, ack => zeropad3D_CP_676_elements(291)); -- 
    cr_3865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(291), ack => type_cast_2066_inst_req_1); -- 
    cr_3956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(291), ack => ptr_deref_2077_load_0_req_1); -- 
    req_4006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(291), ack => array_obj_ref_2097_index_offset_req_1); -- 
    cr_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(291), ack => ptr_deref_2101_store_0_req_1); -- 
    req_3911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(291), ack => addr_of_2073_final_reg_req_1); -- 
    cr_3851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(291), ack => type_cast_2002_inst_req_1); -- 
    rr_3846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(291), ack => type_cast_2002_inst_req_0); -- 
    req_3896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(291), ack => array_obj_ref_2072_index_offset_req_1); -- 
    cr_3975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(291), ack => type_cast_2091_inst_req_1); -- 
    req_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(291), ack => addr_of_2098_final_reg_req_1); -- 
    -- CP-element group 292:  transition  place  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	744 
    -- CP-element group 292:  members (5) 
      -- CP-element group 292: 	 branch_block_stmt_223/if_stmt_1934_else_link/$exit
      -- CP-element group 292: 	 branch_block_stmt_223/if_stmt_1934_else_link/else_choice_transition
      -- CP-element group 292: 	 branch_block_stmt_223/lorx_xlhsx_xfalse769_ifx_xthen786
      -- CP-element group 292: 	 branch_block_stmt_223/lorx_xlhsx_xfalse769_ifx_xthen786_PhiReq/$entry
      -- CP-element group 292: 	 branch_block_stmt_223/lorx_xlhsx_xfalse769_ifx_xthen786_PhiReq/$exit
      -- 
    else_choice_transition_3692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1934_branch_ack_0, ack => zeropad3D_CP_676_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	744 
    -- CP-element group 293: successors 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_Sample/ra
      -- 
    ra_3706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1944_inst_ack_0, ack => zeropad3D_CP_676_elements(293)); -- 
    -- CP-element group 294:  transition  input  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	744 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	297 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_Update/ca
      -- 
    ca_3711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1944_inst_ack_1, ack => zeropad3D_CP_676_elements(294)); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	744 
    -- CP-element group 295: successors 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_Sample/ra
      -- 
    ra_3720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1949_inst_ack_0, ack => zeropad3D_CP_676_elements(295)); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	744 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_Update/ca
      -- 
    ca_3725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1949_inst_ack_1, ack => zeropad3D_CP_676_elements(296)); -- 
    -- CP-element group 297:  join  transition  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	294 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_sample_start_
      -- CP-element group 297: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_Sample/rr
      -- 
    rr_3733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(297), ack => type_cast_1983_inst_req_0); -- 
    zeropad3D_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(294) & zeropad3D_CP_676_elements(296);
      gj_zeropad3D_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_sample_completed_
      -- CP-element group 298: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_Sample/$exit
      -- CP-element group 298: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_Sample/ra
      -- 
    ra_3734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1983_inst_ack_0, ack => zeropad3D_CP_676_elements(298)); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	744 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (16) 
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_update_completed_
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_Update/$exit
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_Update/ca
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_resized_1
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_scaled_1
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_computed_1
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_resize_1/$entry
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_resize_1/$exit
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_resize_1/index_resize_req
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_resize_1/index_resize_ack
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_scale_1/$entry
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_scale_1/$exit
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_scale_1/scale_rename_req
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_index_scale_1/scale_rename_ack
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_final_index_sum_regn_Sample/$entry
      -- CP-element group 299: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_final_index_sum_regn_Sample/req
      -- 
    ca_3739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1983_inst_ack_1, ack => zeropad3D_CP_676_elements(299)); -- 
    req_3764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(299), ack => array_obj_ref_1989_index_offset_req_0); -- 
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	306 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_final_index_sum_regn_sample_complete
      -- CP-element group 300: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_final_index_sum_regn_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_final_index_sum_regn_Sample/ack
      -- 
    ack_3765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1989_index_offset_ack_0, ack => zeropad3D_CP_676_elements(300)); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	744 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (11) 
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_root_address_calculated
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_offset_calculated
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_final_index_sum_regn_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_final_index_sum_regn_Update/ack
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_base_plus_offset/$entry
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_base_plus_offset/$exit
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_base_plus_offset/sum_rename_req
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_base_plus_offset/sum_rename_ack
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_request/$entry
      -- CP-element group 301: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_request/req
      -- 
    ack_3770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1989_index_offset_ack_1, ack => zeropad3D_CP_676_elements(301)); -- 
    req_3779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(301), ack => addr_of_1990_final_reg_req_0); -- 
    -- CP-element group 302:  transition  input  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_sample_completed_
      -- CP-element group 302: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_request/$exit
      -- CP-element group 302: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_request/ack
      -- 
    ack_3780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1990_final_reg_ack_0, ack => zeropad3D_CP_676_elements(302)); -- 
    -- CP-element group 303:  join  fork  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	744 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (28) 
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_word_addrgen/root_register_ack
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/ptr_deref_1993_Split/$entry
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/ptr_deref_1993_Split/$exit
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/ptr_deref_1993_Split/split_req
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/ptr_deref_1993_Split/split_ack
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/word_access_start/$entry
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/word_access_start/word_0/rr
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/word_access_start/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_update_completed_
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_complete/$exit
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_complete/ack
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_base_address_resized
      -- 
    ack_3785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1990_final_reg_ack_1, ack => zeropad3D_CP_676_elements(303)); -- 
    rr_3823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(303), ack => ptr_deref_1993_store_0_req_0); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304:  members (5) 
      -- CP-element group 304: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/$exit
      -- CP-element group 304: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/word_access_start/$exit
      -- CP-element group 304: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/word_access_start/word_0/ra
      -- CP-element group 304: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Sample/word_access_start/word_0/$exit
      -- CP-element group 304: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_sample_completed_
      -- 
    ra_3824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1993_store_0_ack_0, ack => zeropad3D_CP_676_elements(304)); -- 
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	744 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (5) 
      -- CP-element group 305: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Update/word_access_complete/$exit
      -- CP-element group 305: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Update/word_access_complete/word_0/$exit
      -- CP-element group 305: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Update/word_access_complete/word_0/ca
      -- CP-element group 305: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Update/$exit
      -- CP-element group 305: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_update_completed_
      -- 
    ca_3835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1993_store_0_ack_1, ack => zeropad3D_CP_676_elements(305)); -- 
    -- CP-element group 306:  join  transition  place  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	300 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	745 
    -- CP-element group 306:  members (5) 
      -- CP-element group 306: 	 branch_block_stmt_223/ifx_xthen786_ifx_xend855
      -- CP-element group 306: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996__exit__
      -- CP-element group 306: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/$exit
      -- CP-element group 306: 	 branch_block_stmt_223/ifx_xthen786_ifx_xend855_PhiReq/$entry
      -- CP-element group 306: 	 branch_block_stmt_223/ifx_xthen786_ifx_xend855_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(300) & zeropad3D_CP_676_elements(305);
      gj_zeropad3D_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	291 
    -- CP-element group 307: successors 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_Sample/ra
      -- CP-element group 307: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_sample_completed_
      -- 
    ra_3847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2002_inst_ack_0, ack => zeropad3D_CP_676_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	291 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308: 	317 
    -- CP-element group 308:  members (9) 
      -- CP-element group 308: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_Sample/rr
      -- CP-element group 308: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_Update/ca
      -- CP-element group 308: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2002_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_Sample/rr
      -- CP-element group 308: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_Sample/$entry
      -- 
    ca_3852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2002_inst_ack_1, ack => zeropad3D_CP_676_elements(308)); -- 
    rr_3860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(308), ack => type_cast_2066_inst_req_0); -- 
    rr_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(308), ack => type_cast_2091_inst_req_0); -- 
    -- CP-element group 309:  transition  input  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_Sample/ra
      -- CP-element group 309: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_sample_completed_
      -- 
    ra_3861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2066_inst_ack_0, ack => zeropad3D_CP_676_elements(309)); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	291 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (16) 
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_resized_1
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_scaled_1
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_computed_1
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_resize_1/$entry
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_resize_1/$exit
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_Update/ca
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2066_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_final_index_sum_regn_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_final_index_sum_regn_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_scale_1/scale_rename_ack
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_scale_1/scale_rename_req
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_scale_1/$exit
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_scale_1/$entry
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_resize_1/index_resize_ack
      -- CP-element group 310: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_index_resize_1/index_resize_req
      -- 
    ca_3866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2066_inst_ack_1, ack => zeropad3D_CP_676_elements(310)); -- 
    req_3891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(310), ack => array_obj_ref_2072_index_offset_req_0); -- 
    -- CP-element group 311:  transition  input  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	326 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_final_index_sum_regn_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_final_index_sum_regn_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_final_index_sum_regn_sample_complete
      -- 
    ack_3892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2072_index_offset_ack_0, ack => zeropad3D_CP_676_elements(311)); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	291 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (11) 
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_offset_calculated
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_root_address_calculated
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_request/req
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_request/$entry
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_base_plus_offset/sum_rename_ack
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_base_plus_offset/sum_rename_req
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_base_plus_offset/$exit
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_base_plus_offset/$entry
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_final_index_sum_regn_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2072_final_index_sum_regn_Update/$exit
      -- 
    ack_3897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2072_index_offset_ack_1, ack => zeropad3D_CP_676_elements(312)); -- 
    req_3906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(312), ack => addr_of_2073_final_reg_req_0); -- 
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_request/ack
      -- CP-element group 313: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_request/$exit
      -- 
    ack_3907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2073_final_reg_ack_0, ack => zeropad3D_CP_676_elements(313)); -- 
    -- CP-element group 314:  join  fork  transition  input  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	291 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (24) 
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Sample/word_access_start/word_0/rr
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Sample/word_access_start/word_0/$entry
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Sample/word_access_start/$entry
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Sample/$entry
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_word_addrgen/root_register_ack
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_word_addrgen/root_register_req
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_word_addrgen/$exit
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_word_addrgen/$entry
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_base_plus_offset/sum_rename_ack
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_base_plus_offset/sum_rename_req
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_base_plus_offset/$exit
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_base_plus_offset/$entry
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_base_addr_resize/base_resize_ack
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_base_addr_resize/base_resize_req
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_base_addr_resize/$exit
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_base_addr_resize/$entry
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_base_address_resized
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_root_address_calculated
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_word_address_calculated
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_base_address_calculated
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_sample_start_
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_complete/ack
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_complete/$exit
      -- CP-element group 314: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2073_update_completed_
      -- 
    ack_3912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2073_final_reg_ack_1, ack => zeropad3D_CP_676_elements(314)); -- 
    rr_3945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(314), ack => ptr_deref_2077_load_0_req_0); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (5) 
      -- CP-element group 315: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Sample/word_access_start/word_0/ra
      -- CP-element group 315: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Sample/word_access_start/word_0/$exit
      -- CP-element group 315: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Sample/word_access_start/$exit
      -- CP-element group 315: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_sample_completed_
      -- 
    ra_3946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2077_load_0_ack_0, ack => zeropad3D_CP_676_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	291 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	323 
    -- CP-element group 316:  members (9) 
      -- CP-element group 316: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/ptr_deref_2077_Merge/$entry
      -- CP-element group 316: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/ptr_deref_2077_Merge/$exit
      -- CP-element group 316: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/ptr_deref_2077_Merge/merge_req
      -- CP-element group 316: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/ptr_deref_2077_Merge/merge_ack
      -- CP-element group 316: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/word_access_complete/$exit
      -- CP-element group 316: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/word_access_complete/word_0/$exit
      -- CP-element group 316: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2077_Update/word_access_complete/word_0/ca
      -- 
    ca_3957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2077_load_0_ack_1, ack => zeropad3D_CP_676_elements(316)); -- 
    -- CP-element group 317:  transition  input  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	308 
    -- CP-element group 317: successors 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_sample_completed_
      -- CP-element group 317: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_Sample/ra
      -- CP-element group 317: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_Sample/$exit
      -- 
    ra_3971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2091_inst_ack_0, ack => zeropad3D_CP_676_elements(317)); -- 
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	291 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (16) 
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_update_completed_
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_final_index_sum_regn_Sample/req
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_final_index_sum_regn_Sample/$entry
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_scale_1/scale_rename_ack
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_scale_1/scale_rename_req
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_scale_1/$exit
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_scale_1/$entry
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_resize_1/index_resize_ack
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_resize_1/index_resize_req
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_resize_1/$exit
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_resize_1/$entry
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_computed_1
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_scaled_1
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_index_resized_1
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_Update/ca
      -- CP-element group 318: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/type_cast_2091_Update/$exit
      -- 
    ca_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2091_inst_ack_1, ack => zeropad3D_CP_676_elements(318)); -- 
    req_4001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(318), ack => array_obj_ref_2097_index_offset_req_0); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	326 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_final_index_sum_regn_Sample/ack
      -- CP-element group 319: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_final_index_sum_regn_Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_final_index_sum_regn_sample_complete
      -- 
    ack_4002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2097_index_offset_ack_0, ack => zeropad3D_CP_676_elements(319)); -- 
    -- CP-element group 320:  transition  input  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	291 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (11) 
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_final_index_sum_regn_Update/ack
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_base_plus_offset/$entry
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_base_plus_offset/$exit
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_base_plus_offset/sum_rename_req
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_base_plus_offset/sum_rename_ack
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_request/$entry
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_request/req
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_final_index_sum_regn_Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_offset_calculated
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/array_obj_ref_2097_root_address_calculated
      -- CP-element group 320: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_sample_start_
      -- 
    ack_4007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2097_index_offset_ack_1, ack => zeropad3D_CP_676_elements(320)); -- 
    req_4016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(320), ack => addr_of_2098_final_reg_req_0); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_request/$exit
      -- CP-element group 321: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_request/ack
      -- CP-element group 321: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_sample_completed_
      -- 
    ack_4017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2098_final_reg_ack_0, ack => zeropad3D_CP_676_elements(321)); -- 
    -- CP-element group 322:  fork  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	291 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (19) 
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_base_plus_offset/$entry
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_base_plus_offset/$exit
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_base_plus_offset/sum_rename_req
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_base_plus_offset/sum_rename_ack
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_complete/$exit
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_word_addrgen/$entry
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_word_addrgen/$exit
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_base_addr_resize/base_resize_ack
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_base_addr_resize/base_resize_req
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_base_addr_resize/$exit
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_word_addrgen/root_register_ack
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_base_addr_resize/$entry
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_base_address_resized
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_root_address_calculated
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_word_address_calculated
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_base_address_calculated
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_update_completed_
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_word_addrgen/root_register_req
      -- CP-element group 322: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/addr_of_2098_complete/ack
      -- 
    ack_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2098_final_reg_ack_1, ack => zeropad3D_CP_676_elements(322)); -- 
    -- CP-element group 323:  join  transition  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	316 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (9) 
      -- CP-element group 323: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/ptr_deref_2101_Split/split_ack
      -- CP-element group 323: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/ptr_deref_2101_Split/$entry
      -- CP-element group 323: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/ptr_deref_2101_Split/$exit
      -- CP-element group 323: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/ptr_deref_2101_Split/split_req
      -- CP-element group 323: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/$entry
      -- CP-element group 323: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/word_access_start/word_0/rr
      -- CP-element group 323: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_sample_start_
      -- CP-element group 323: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/word_access_start/$entry
      -- CP-element group 323: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/word_access_start/word_0/$entry
      -- 
    rr_4060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(323), ack => ptr_deref_2101_store_0_req_0); -- 
    zeropad3D_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(316) & zeropad3D_CP_676_elements(322);
      gj_zeropad3D_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324:  members (5) 
      -- CP-element group 324: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/word_access_start/word_0/ra
      -- CP-element group 324: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/word_access_start/word_0/$exit
      -- CP-element group 324: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_sample_completed_
      -- CP-element group 324: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Sample/word_access_start/$exit
      -- 
    ra_4061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2101_store_0_ack_0, ack => zeropad3D_CP_676_elements(324)); -- 
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	291 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (5) 
      -- CP-element group 325: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Update/word_access_complete/word_0/ca
      -- CP-element group 325: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Update/word_access_complete/word_0/$exit
      -- CP-element group 325: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Update/word_access_complete/$exit
      -- CP-element group 325: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/ptr_deref_2101_update_completed_
      -- 
    ca_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2101_store_0_ack_1, ack => zeropad3D_CP_676_elements(325)); -- 
    -- CP-element group 326:  join  transition  place  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	311 
    -- CP-element group 326: 	319 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	745 
    -- CP-element group 326:  members (5) 
      -- CP-element group 326: 	 branch_block_stmt_223/ifx_xelse807_ifx_xend855
      -- CP-element group 326: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103__exit__
      -- CP-element group 326: 	 branch_block_stmt_223/assign_stmt_2003_to_assign_stmt_2103/$exit
      -- CP-element group 326: 	 branch_block_stmt_223/ifx_xelse807_ifx_xend855_PhiReq/$entry
      -- CP-element group 326: 	 branch_block_stmt_223/ifx_xelse807_ifx_xend855_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(311) & zeropad3D_CP_676_elements(319) & zeropad3D_CP_676_elements(325);
      gj_zeropad3D_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	745 
    -- CP-element group 327: successors 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_Sample/ra
      -- 
    ra_4084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2109_inst_ack_0, ack => zeropad3D_CP_676_elements(327)); -- 
    -- CP-element group 328:  branch  transition  place  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	745 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328: 	330 
    -- CP-element group 328:  members (13) 
      -- CP-element group 328: 	 branch_block_stmt_223/if_stmt_2124__entry__
      -- CP-element group 328: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123__exit__
      -- CP-element group 328: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_223/if_stmt_2124_if_link/$entry
      -- CP-element group 328: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/$exit
      -- CP-element group 328: 	 branch_block_stmt_223/if_stmt_2124_else_link/$entry
      -- CP-element group 328: 	 branch_block_stmt_223/if_stmt_2124_eval_test/branch_req
      -- CP-element group 328: 	 branch_block_stmt_223/if_stmt_2124_eval_test/$exit
      -- CP-element group 328: 	 branch_block_stmt_223/if_stmt_2124_eval_test/$entry
      -- CP-element group 328: 	 branch_block_stmt_223/R_cmp863_2125_place
      -- CP-element group 328: 	 branch_block_stmt_223/if_stmt_2124_dead_link/$entry
      -- CP-element group 328: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_Update/ca
      -- CP-element group 328: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_Update/$exit
      -- 
    ca_4089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2109_inst_ack_1, ack => zeropad3D_CP_676_elements(328)); -- 
    branch_req_4097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(328), ack => if_stmt_2124_branch_req_0); -- 
    -- CP-element group 329:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	754 
    -- CP-element group 329: 	755 
    -- CP-element group 329: 	757 
    -- CP-element group 329: 	758 
    -- CP-element group 329: 	760 
    -- CP-element group 329: 	761 
    -- CP-element group 329:  members (40) 
      -- CP-element group 329: 	 branch_block_stmt_223/assign_stmt_2136__entry__
      -- CP-element group 329: 	 branch_block_stmt_223/assign_stmt_2136__exit__
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906
      -- CP-element group 329: 	 branch_block_stmt_223/merge_stmt_2130__exit__
      -- CP-element group 329: 	 branch_block_stmt_223/if_stmt_2124_if_link/$exit
      -- CP-element group 329: 	 branch_block_stmt_223/assign_stmt_2136/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/assign_stmt_2136/$exit
      -- CP-element group 329: 	 branch_block_stmt_223/if_stmt_2124_if_link/if_choice_transition
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xend855_ifx_xthen865
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xend855_ifx_xthen865_PhiReq/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xend855_ifx_xthen865_PhiReq/$exit
      -- CP-element group 329: 	 branch_block_stmt_223/merge_stmt_2130_PhiReqMerge
      -- CP-element group 329: 	 branch_block_stmt_223/merge_stmt_2130_PhiAck/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/merge_stmt_2130_PhiAck/$exit
      -- CP-element group 329: 	 branch_block_stmt_223/merge_stmt_2130_PhiAck/dummy
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/SplitProtocol/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/SplitProtocol/Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/SplitProtocol/Sample/rr
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/SplitProtocol/Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/SplitProtocol/Update/cr
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/rr
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/cr
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/SplitProtocol/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/SplitProtocol/Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/SplitProtocol/Sample/rr
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/SplitProtocol/Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2124_branch_ack_1, ack => zeropad3D_CP_676_elements(329)); -- 
    rr_7981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(329), ack => type_cast_2193_inst_req_0); -- 
    cr_7986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(329), ack => type_cast_2193_inst_req_1); -- 
    rr_8004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(329), ack => type_cast_2197_inst_req_0); -- 
    cr_8009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(329), ack => type_cast_2197_inst_req_1); -- 
    rr_8027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(329), ack => type_cast_2205_inst_req_0); -- 
    cr_8032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(329), ack => type_cast_2205_inst_req_1); -- 
    -- CP-element group 330:  fork  transition  place  input  output  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	328 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330: 	332 
    -- CP-element group 330: 	334 
    -- CP-element group 330: 	336 
    -- CP-element group 330:  members (24) 
      -- CP-element group 330: 	 branch_block_stmt_223/merge_stmt_2138__exit__
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179__entry__
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/$entry
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_sample_start_
      -- CP-element group 330: 	 branch_block_stmt_223/if_stmt_2124_else_link/$exit
      -- CP-element group 330: 	 branch_block_stmt_223/if_stmt_2124_else_link/else_choice_transition
      -- CP-element group 330: 	 branch_block_stmt_223/ifx_xend855_ifx_xelse870
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_update_start_
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_Sample/$entry
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_Sample/rr
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_Update/cr
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_update_start_
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_Update/cr
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_update_start_
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_Update/cr
      -- CP-element group 330: 	 branch_block_stmt_223/ifx_xend855_ifx_xelse870_PhiReq/$entry
      -- CP-element group 330: 	 branch_block_stmt_223/ifx_xend855_ifx_xelse870_PhiReq/$exit
      -- CP-element group 330: 	 branch_block_stmt_223/merge_stmt_2138_PhiReqMerge
      -- CP-element group 330: 	 branch_block_stmt_223/merge_stmt_2138_PhiAck/$entry
      -- CP-element group 330: 	 branch_block_stmt_223/merge_stmt_2138_PhiAck/$exit
      -- CP-element group 330: 	 branch_block_stmt_223/merge_stmt_2138_PhiAck/dummy
      -- 
    else_choice_transition_4106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2124_branch_ack_0, ack => zeropad3D_CP_676_elements(330)); -- 
    rr_4122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(330), ack => type_cast_2148_inst_req_0); -- 
    cr_4127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(330), ack => type_cast_2148_inst_req_1); -- 
    cr_4141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(330), ack => type_cast_2157_inst_req_1); -- 
    cr_4155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(330), ack => type_cast_2173_inst_req_1); -- 
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_Sample/ra
      -- 
    ra_4123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2148_inst_ack_0, ack => zeropad3D_CP_676_elements(331)); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2148_Update/ca
      -- CP-element group 332: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_Sample/rr
      -- 
    ca_4128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2148_inst_ack_1, ack => zeropad3D_CP_676_elements(332)); -- 
    rr_4136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(332), ack => type_cast_2157_inst_req_0); -- 
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_Sample/ra
      -- 
    ra_4137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2157_inst_ack_0, ack => zeropad3D_CP_676_elements(333)); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	330 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2157_Update/ca
      -- CP-element group 334: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_Sample/rr
      -- 
    ca_4142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2157_inst_ack_1, ack => zeropad3D_CP_676_elements(334)); -- 
    rr_4150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(334), ack => type_cast_2173_inst_req_0); -- 
    -- CP-element group 335:  transition  input  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_Sample/ra
      -- 
    ra_4151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2173_inst_ack_0, ack => zeropad3D_CP_676_elements(335)); -- 
    -- CP-element group 336:  branch  transition  place  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	330 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336: 	338 
    -- CP-element group 336:  members (13) 
      -- CP-element group 336: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179__exit__
      -- CP-element group 336: 	 branch_block_stmt_223/if_stmt_2180__entry__
      -- CP-element group 336: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/$exit
      -- CP-element group 336: 	 branch_block_stmt_223/R_cmp897_2181_place
      -- CP-element group 336: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_223/assign_stmt_2144_to_assign_stmt_2179/type_cast_2173_Update/ca
      -- CP-element group 336: 	 branch_block_stmt_223/if_stmt_2180_dead_link/$entry
      -- CP-element group 336: 	 branch_block_stmt_223/if_stmt_2180_eval_test/$entry
      -- CP-element group 336: 	 branch_block_stmt_223/if_stmt_2180_eval_test/$exit
      -- CP-element group 336: 	 branch_block_stmt_223/if_stmt_2180_eval_test/branch_req
      -- CP-element group 336: 	 branch_block_stmt_223/if_stmt_2180_if_link/$entry
      -- CP-element group 336: 	 branch_block_stmt_223/if_stmt_2180_else_link/$entry
      -- 
    ca_4156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2173_inst_ack_1, ack => zeropad3D_CP_676_elements(336)); -- 
    branch_req_4164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(336), ack => if_stmt_2180_branch_req_0); -- 
    -- CP-element group 337:  fork  transition  place  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	339 
    -- CP-element group 337: 	340 
    -- CP-element group 337: 	342 
    -- CP-element group 337:  members (27) 
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259__entry__
      -- CP-element group 337: 	 branch_block_stmt_223/merge_stmt_2208__exit__
      -- CP-element group 337: 	 branch_block_stmt_223/ifx_xelse870_whilex_xend907
      -- CP-element group 337: 	 branch_block_stmt_223/if_stmt_2180_if_link/$exit
      -- CP-element group 337: 	 branch_block_stmt_223/if_stmt_2180_if_link/if_choice_transition
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/$entry
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_update_start_
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_word_address_calculated
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_root_address_calculated
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Sample/word_access_start/$entry
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Sample/word_access_start/word_0/$entry
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Sample/word_access_start/word_0/rr
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/word_access_complete/$entry
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/word_access_complete/word_0/$entry
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/word_access_complete/word_0/cr
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_update_start_
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_Update/cr
      -- CP-element group 337: 	 branch_block_stmt_223/ifx_xelse870_whilex_xend907_PhiReq/$entry
      -- CP-element group 337: 	 branch_block_stmt_223/ifx_xelse870_whilex_xend907_PhiReq/$exit
      -- CP-element group 337: 	 branch_block_stmt_223/merge_stmt_2208_PhiReqMerge
      -- CP-element group 337: 	 branch_block_stmt_223/merge_stmt_2208_PhiAck/$entry
      -- CP-element group 337: 	 branch_block_stmt_223/merge_stmt_2208_PhiAck/$exit
      -- CP-element group 337: 	 branch_block_stmt_223/merge_stmt_2208_PhiAck/dummy
      -- 
    if_choice_transition_4169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2180_branch_ack_1, ack => zeropad3D_CP_676_elements(337)); -- 
    rr_4194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(337), ack => LOAD_pad_2216_load_0_req_0); -- 
    cr_4205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(337), ack => LOAD_pad_2216_load_0_req_1); -- 
    cr_4224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(337), ack => type_cast_2220_inst_req_1); -- 
    -- CP-element group 338:  fork  transition  place  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	336 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	746 
    -- CP-element group 338: 	747 
    -- CP-element group 338: 	748 
    -- CP-element group 338: 	750 
    -- CP-element group 338: 	751 
    -- CP-element group 338:  members (22) 
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906
      -- CP-element group 338: 	 branch_block_stmt_223/if_stmt_2180_else_link/$exit
      -- CP-element group 338: 	 branch_block_stmt_223/if_stmt_2180_else_link/else_choice_transition
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2187/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/rr
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/cr
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/SplitProtocol/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/SplitProtocol/Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/SplitProtocol/Sample/rr
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/SplitProtocol/Update/$entry
      -- CP-element group 338: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2180_branch_ack_0, ack => zeropad3D_CP_676_elements(338)); -- 
    rr_7932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(338), ack => type_cast_2199_inst_req_0); -- 
    cr_7937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(338), ack => type_cast_2199_inst_req_1); -- 
    rr_7955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(338), ack => type_cast_2203_inst_req_0); -- 
    cr_7960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(338), ack => type_cast_2203_inst_req_1); -- 
    -- CP-element group 339:  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	337 
    -- CP-element group 339: successors 
    -- CP-element group 339:  members (5) 
      -- CP-element group 339: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Sample/word_access_start/$exit
      -- CP-element group 339: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Sample/word_access_start/word_0/$exit
      -- CP-element group 339: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Sample/word_access_start/word_0/ra
      -- 
    ra_4195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2216_load_0_ack_0, ack => zeropad3D_CP_676_elements(339)); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	337 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (12) 
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/word_access_complete/$exit
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/word_access_complete/word_0/$exit
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/word_access_complete/word_0/ca
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/LOAD_pad_2216_Merge/$entry
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/LOAD_pad_2216_Merge/$exit
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/LOAD_pad_2216_Merge/merge_req
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/LOAD_pad_2216_Update/LOAD_pad_2216_Merge/merge_ack
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_Sample/rr
      -- 
    ca_4206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2216_load_0_ack_1, ack => zeropad3D_CP_676_elements(340)); -- 
    rr_4219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(340), ack => type_cast_2220_inst_req_0); -- 
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_Sample/ra
      -- 
    ra_4220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2220_inst_ack_0, ack => zeropad3D_CP_676_elements(341)); -- 
    -- CP-element group 342:  fork  transition  place  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	337 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	779 
    -- CP-element group 342: 	780 
    -- CP-element group 342: 	781 
    -- CP-element group 342: 	783 
    -- CP-element group 342:  members (19) 
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967
      -- CP-element group 342: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259__exit__
      -- CP-element group 342: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/$exit
      -- CP-element group 342: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_223/assign_stmt_2214_to_assign_stmt_2259/type_cast_2220_Update/ca
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/$entry
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2262/$entry
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/$entry
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/$entry
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/$entry
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/$entry
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/$entry
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Sample/rr
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Update/$entry
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Update/cr
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2275/$entry
      -- CP-element group 342: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/$entry
      -- 
    ca_4225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2220_inst_ack_1, ack => zeropad3D_CP_676_elements(342)); -- 
    rr_8148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(342), ack => type_cast_2272_inst_req_0); -- 
    cr_8153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(342), ack => type_cast_2272_inst_req_1); -- 
    -- CP-element group 343:  transition  input  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	789 
    -- CP-element group 343: successors 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_Sample/ra
      -- 
    ra_4237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2286_inst_ack_0, ack => zeropad3D_CP_676_elements(343)); -- 
    -- CP-element group 344:  branch  transition  place  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	789 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344: 	346 
    -- CP-element group 344:  members (13) 
      -- CP-element group 344: 	 branch_block_stmt_223/if_stmt_2313__entry__
      -- CP-element group 344: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312__exit__
      -- CP-element group 344: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/$exit
      -- CP-element group 344: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_Update/ca
      -- CP-element group 344: 	 branch_block_stmt_223/if_stmt_2313_dead_link/$entry
      -- CP-element group 344: 	 branch_block_stmt_223/if_stmt_2313_eval_test/$entry
      -- CP-element group 344: 	 branch_block_stmt_223/if_stmt_2313_eval_test/$exit
      -- CP-element group 344: 	 branch_block_stmt_223/if_stmt_2313_eval_test/branch_req
      -- CP-element group 344: 	 branch_block_stmt_223/R_orx_xcond1856_2314_place
      -- CP-element group 344: 	 branch_block_stmt_223/if_stmt_2313_if_link/$entry
      -- CP-element group 344: 	 branch_block_stmt_223/if_stmt_2313_else_link/$entry
      -- 
    ca_4242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2286_inst_ack_1, ack => zeropad3D_CP_676_elements(344)); -- 
    branch_req_4250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(344), ack => if_stmt_2313_branch_req_0); -- 
    -- CP-element group 345:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	347 
    -- CP-element group 345: 	348 
    -- CP-element group 345:  members (18) 
      -- CP-element group 345: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349__entry__
      -- CP-element group 345: 	 branch_block_stmt_223/merge_stmt_2319__exit__
      -- CP-element group 345: 	 branch_block_stmt_223/if_stmt_2313_if_link/$exit
      -- CP-element group 345: 	 branch_block_stmt_223/if_stmt_2313_if_link/if_choice_transition
      -- CP-element group 345: 	 branch_block_stmt_223/whilex_xbody967_lorx_xlhsx_xfalse986
      -- CP-element group 345: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/$entry
      -- CP-element group 345: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_sample_start_
      -- CP-element group 345: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_update_start_
      -- CP-element group 345: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_Sample/rr
      -- CP-element group 345: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_Update/cr
      -- CP-element group 345: 	 branch_block_stmt_223/whilex_xbody967_lorx_xlhsx_xfalse986_PhiReq/$entry
      -- CP-element group 345: 	 branch_block_stmt_223/whilex_xbody967_lorx_xlhsx_xfalse986_PhiReq/$exit
      -- CP-element group 345: 	 branch_block_stmt_223/merge_stmt_2319_PhiReqMerge
      -- CP-element group 345: 	 branch_block_stmt_223/merge_stmt_2319_PhiAck/$entry
      -- CP-element group 345: 	 branch_block_stmt_223/merge_stmt_2319_PhiAck/$exit
      -- CP-element group 345: 	 branch_block_stmt_223/merge_stmt_2319_PhiAck/dummy
      -- 
    if_choice_transition_4255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2313_branch_ack_1, ack => zeropad3D_CP_676_elements(345)); -- 
    rr_4272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(345), ack => type_cast_2323_inst_req_0); -- 
    cr_4277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(345), ack => type_cast_2323_inst_req_1); -- 
    -- CP-element group 346:  transition  place  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	344 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	790 
    -- CP-element group 346:  members (5) 
      -- CP-element group 346: 	 branch_block_stmt_223/if_stmt_2313_else_link/$exit
      -- CP-element group 346: 	 branch_block_stmt_223/if_stmt_2313_else_link/else_choice_transition
      -- CP-element group 346: 	 branch_block_stmt_223/whilex_xbody967_ifx_xthen1004
      -- CP-element group 346: 	 branch_block_stmt_223/whilex_xbody967_ifx_xthen1004_PhiReq/$entry
      -- CP-element group 346: 	 branch_block_stmt_223/whilex_xbody967_ifx_xthen1004_PhiReq/$exit
      -- 
    else_choice_transition_4259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2313_branch_ack_0, ack => zeropad3D_CP_676_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_Sample/ra
      -- 
    ra_4273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2323_inst_ack_0, ack => zeropad3D_CP_676_elements(347)); -- 
    -- CP-element group 348:  branch  transition  place  input  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	345 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348: 	350 
    -- CP-element group 348:  members (13) 
      -- CP-element group 348: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349__exit__
      -- CP-element group 348: 	 branch_block_stmt_223/if_stmt_2350__entry__
      -- CP-element group 348: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/$exit
      -- CP-element group 348: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_223/assign_stmt_2324_to_assign_stmt_2349/type_cast_2323_Update/ca
      -- CP-element group 348: 	 branch_block_stmt_223/if_stmt_2350_dead_link/$entry
      -- CP-element group 348: 	 branch_block_stmt_223/if_stmt_2350_eval_test/$entry
      -- CP-element group 348: 	 branch_block_stmt_223/if_stmt_2350_eval_test/$exit
      -- CP-element group 348: 	 branch_block_stmt_223/if_stmt_2350_eval_test/branch_req
      -- CP-element group 348: 	 branch_block_stmt_223/R_orx_xcond1857_2351_place
      -- CP-element group 348: 	 branch_block_stmt_223/if_stmt_2350_if_link/$entry
      -- CP-element group 348: 	 branch_block_stmt_223/if_stmt_2350_else_link/$entry
      -- 
    ca_4278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2323_inst_ack_1, ack => zeropad3D_CP_676_elements(348)); -- 
    branch_req_4286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(348), ack => if_stmt_2350_branch_req_0); -- 
    -- CP-element group 349:  fork  transition  place  input  output  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	365 
    -- CP-element group 349: 	366 
    -- CP-element group 349: 	368 
    -- CP-element group 349: 	370 
    -- CP-element group 349: 	372 
    -- CP-element group 349: 	374 
    -- CP-element group 349: 	376 
    -- CP-element group 349: 	378 
    -- CP-element group 349: 	380 
    -- CP-element group 349: 	383 
    -- CP-element group 349:  members (46) 
      -- CP-element group 349: 	 branch_block_stmt_223/merge_stmt_2414__exit__
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519__entry__
      -- CP-element group 349: 	 branch_block_stmt_223/if_stmt_2350_if_link/$exit
      -- CP-element group 349: 	 branch_block_stmt_223/if_stmt_2350_if_link/if_choice_transition
      -- CP-element group 349: 	 branch_block_stmt_223/lorx_xlhsx_xfalse986_ifx_xelse1025
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_sample_start_
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_update_start_
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_Sample/rr
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_Update/cr
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_update_start_
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_Update/cr
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_update_start_
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_final_index_sum_regn_update_start
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_final_index_sum_regn_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_final_index_sum_regn_Update/req
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_complete/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_complete/req
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_update_start_
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/word_access_complete/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/word_access_complete/word_0/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/word_access_complete/word_0/cr
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_update_start_
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_Update/cr
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_update_start_
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_final_index_sum_regn_update_start
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_final_index_sum_regn_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_final_index_sum_regn_Update/req
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_complete/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_complete/req
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_update_start_
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Update/word_access_complete/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Update/word_access_complete/word_0/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Update/word_access_complete/word_0/cr
      -- CP-element group 349: 	 branch_block_stmt_223/lorx_xlhsx_xfalse986_ifx_xelse1025_PhiReq/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/lorx_xlhsx_xfalse986_ifx_xelse1025_PhiReq/$exit
      -- CP-element group 349: 	 branch_block_stmt_223/merge_stmt_2414_PhiReqMerge
      -- CP-element group 349: 	 branch_block_stmt_223/merge_stmt_2414_PhiAck/$entry
      -- CP-element group 349: 	 branch_block_stmt_223/merge_stmt_2414_PhiAck/$exit
      -- CP-element group 349: 	 branch_block_stmt_223/merge_stmt_2414_PhiAck/dummy
      -- 
    if_choice_transition_4291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2350_branch_ack_1, ack => zeropad3D_CP_676_elements(349)); -- 
    rr_4449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => type_cast_2418_inst_req_0); -- 
    cr_4454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => type_cast_2418_inst_req_1); -- 
    cr_4468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => type_cast_2482_inst_req_1); -- 
    req_4499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => array_obj_ref_2488_index_offset_req_1); -- 
    req_4514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => addr_of_2489_final_reg_req_1); -- 
    cr_4559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => ptr_deref_2493_load_0_req_1); -- 
    cr_4578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => type_cast_2507_inst_req_1); -- 
    req_4609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => array_obj_ref_2513_index_offset_req_1); -- 
    req_4624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => addr_of_2514_final_reg_req_1); -- 
    cr_4674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(349), ack => ptr_deref_2517_store_0_req_1); -- 
    -- CP-element group 350:  transition  place  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	348 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	790 
    -- CP-element group 350:  members (5) 
      -- CP-element group 350: 	 branch_block_stmt_223/if_stmt_2350_else_link/$exit
      -- CP-element group 350: 	 branch_block_stmt_223/if_stmt_2350_else_link/else_choice_transition
      -- CP-element group 350: 	 branch_block_stmt_223/lorx_xlhsx_xfalse986_ifx_xthen1004
      -- CP-element group 350: 	 branch_block_stmt_223/lorx_xlhsx_xfalse986_ifx_xthen1004_PhiReq/$entry
      -- CP-element group 350: 	 branch_block_stmt_223/lorx_xlhsx_xfalse986_ifx_xthen1004_PhiReq/$exit
      -- 
    else_choice_transition_4295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2350_branch_ack_0, ack => zeropad3D_CP_676_elements(350)); -- 
    -- CP-element group 351:  transition  input  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	790 
    -- CP-element group 351: successors 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_sample_completed_
      -- CP-element group 351: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_Sample/ra
      -- 
    ra_4309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2360_inst_ack_0, ack => zeropad3D_CP_676_elements(351)); -- 
    -- CP-element group 352:  transition  input  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	790 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	355 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_update_completed_
      -- CP-element group 352: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_Update/ca
      -- 
    ca_4314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2360_inst_ack_1, ack => zeropad3D_CP_676_elements(352)); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	790 
    -- CP-element group 353: successors 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_sample_completed_
      -- CP-element group 353: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_Sample/$exit
      -- CP-element group 353: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_Sample/ra
      -- 
    ra_4323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2365_inst_ack_0, ack => zeropad3D_CP_676_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	790 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_update_completed_
      -- CP-element group 354: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_Update/$exit
      -- CP-element group 354: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_Update/ca
      -- 
    ca_4328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2365_inst_ack_1, ack => zeropad3D_CP_676_elements(354)); -- 
    -- CP-element group 355:  join  transition  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	352 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_Sample/rr
      -- 
    rr_4336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(355), ack => type_cast_2399_inst_req_0); -- 
    zeropad3D_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(352) & zeropad3D_CP_676_elements(354);
      gj_zeropad3D_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_Sample/ra
      -- 
    ra_4337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2399_inst_ack_0, ack => zeropad3D_CP_676_elements(356)); -- 
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	790 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (16) 
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_Update/ca
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_resized_1
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_scaled_1
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_computed_1
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_resize_1/$entry
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_resize_1/$exit
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_resize_1/index_resize_req
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_resize_1/index_resize_ack
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_scale_1/$entry
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_scale_1/$exit
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_scale_1/scale_rename_req
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_index_scale_1/scale_rename_ack
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_final_index_sum_regn_Sample/$entry
      -- CP-element group 357: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_final_index_sum_regn_Sample/req
      -- 
    ca_4342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2399_inst_ack_1, ack => zeropad3D_CP_676_elements(357)); -- 
    req_4367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(357), ack => array_obj_ref_2405_index_offset_req_0); -- 
    -- CP-element group 358:  transition  input  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	364 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_final_index_sum_regn_sample_complete
      -- CP-element group 358: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_final_index_sum_regn_Sample/$exit
      -- CP-element group 358: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_final_index_sum_regn_Sample/ack
      -- 
    ack_4368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2405_index_offset_ack_0, ack => zeropad3D_CP_676_elements(358)); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	790 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (11) 
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_sample_start_
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_root_address_calculated
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_offset_calculated
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_final_index_sum_regn_Update/$exit
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_final_index_sum_regn_Update/ack
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_base_plus_offset/$entry
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_base_plus_offset/$exit
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_base_plus_offset/sum_rename_req
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_base_plus_offset/sum_rename_ack
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_request/$entry
      -- CP-element group 359: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_request/req
      -- 
    ack_4373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2405_index_offset_ack_1, ack => zeropad3D_CP_676_elements(359)); -- 
    req_4382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(359), ack => addr_of_2406_final_reg_req_0); -- 
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_sample_completed_
      -- CP-element group 360: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_request/$exit
      -- CP-element group 360: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_request/ack
      -- 
    ack_4383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2406_final_reg_ack_0, ack => zeropad3D_CP_676_elements(360)); -- 
    -- CP-element group 361:  join  fork  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	790 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (28) 
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_update_completed_
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_complete/$exit
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_complete/ack
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_sample_start_
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_base_address_calculated
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_word_address_calculated
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_root_address_calculated
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_base_address_resized
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_base_addr_resize/$entry
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_base_addr_resize/$exit
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_base_addr_resize/base_resize_req
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_base_addr_resize/base_resize_ack
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_base_plus_offset/$entry
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_base_plus_offset/$exit
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_base_plus_offset/sum_rename_req
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_base_plus_offset/sum_rename_ack
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_word_addrgen/$entry
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_word_addrgen/$exit
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_word_addrgen/root_register_req
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_word_addrgen/root_register_ack
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/$entry
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/ptr_deref_2409_Split/$entry
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/ptr_deref_2409_Split/$exit
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/ptr_deref_2409_Split/split_req
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/ptr_deref_2409_Split/split_ack
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/word_access_start/$entry
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/word_access_start/word_0/$entry
      -- CP-element group 361: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/word_access_start/word_0/rr
      -- 
    ack_4388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2406_final_reg_ack_1, ack => zeropad3D_CP_676_elements(361)); -- 
    rr_4426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(361), ack => ptr_deref_2409_store_0_req_0); -- 
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362:  members (5) 
      -- CP-element group 362: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_sample_completed_
      -- CP-element group 362: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/word_access_start/$exit
      -- CP-element group 362: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/word_access_start/word_0/$exit
      -- CP-element group 362: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Sample/word_access_start/word_0/ra
      -- 
    ra_4427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2409_store_0_ack_0, ack => zeropad3D_CP_676_elements(362)); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	790 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (5) 
      -- CP-element group 363: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_update_completed_
      -- CP-element group 363: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Update/word_access_complete/$exit
      -- CP-element group 363: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Update/word_access_complete/word_0/$exit
      -- CP-element group 363: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Update/word_access_complete/word_0/ca
      -- 
    ca_4438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2409_store_0_ack_1, ack => zeropad3D_CP_676_elements(363)); -- 
    -- CP-element group 364:  join  transition  place  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	358 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	791 
    -- CP-element group 364:  members (5) 
      -- CP-element group 364: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412__exit__
      -- CP-element group 364: 	 branch_block_stmt_223/ifx_xthen1004_ifx_xend1073
      -- CP-element group 364: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/$exit
      -- CP-element group 364: 	 branch_block_stmt_223/ifx_xthen1004_ifx_xend1073_PhiReq/$entry
      -- CP-element group 364: 	 branch_block_stmt_223/ifx_xthen1004_ifx_xend1073_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(358) & zeropad3D_CP_676_elements(363);
      gj_zeropad3D_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  transition  input  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	349 
    -- CP-element group 365: successors 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_Sample/ra
      -- 
    ra_4450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2418_inst_ack_0, ack => zeropad3D_CP_676_elements(365)); -- 
    -- CP-element group 366:  fork  transition  input  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	349 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366: 	375 
    -- CP-element group 366:  members (9) 
      -- CP-element group 366: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2418_Update/ca
      -- CP-element group 366: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_Sample/rr
      -- CP-element group 366: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_Sample/rr
      -- 
    ca_4455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2418_inst_ack_1, ack => zeropad3D_CP_676_elements(366)); -- 
    rr_4463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(366), ack => type_cast_2482_inst_req_0); -- 
    rr_4573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(366), ack => type_cast_2507_inst_req_0); -- 
    -- CP-element group 367:  transition  input  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_Sample/ra
      -- 
    ra_4464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2482_inst_ack_0, ack => zeropad3D_CP_676_elements(367)); -- 
    -- CP-element group 368:  transition  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	349 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (16) 
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2482_Update/ca
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_resized_1
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_scaled_1
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_computed_1
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_resize_1/$entry
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_resize_1/$exit
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_resize_1/index_resize_req
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_resize_1/index_resize_ack
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_scale_1/$entry
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_scale_1/$exit
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_scale_1/scale_rename_req
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_index_scale_1/scale_rename_ack
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_final_index_sum_regn_Sample/$entry
      -- CP-element group 368: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_final_index_sum_regn_Sample/req
      -- 
    ca_4469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2482_inst_ack_1, ack => zeropad3D_CP_676_elements(368)); -- 
    req_4494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(368), ack => array_obj_ref_2488_index_offset_req_0); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	384 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_final_index_sum_regn_sample_complete
      -- CP-element group 369: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_final_index_sum_regn_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_final_index_sum_regn_Sample/ack
      -- 
    ack_4495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2488_index_offset_ack_0, ack => zeropad3D_CP_676_elements(369)); -- 
    -- CP-element group 370:  transition  input  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	349 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (11) 
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_sample_start_
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_root_address_calculated
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_offset_calculated
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_final_index_sum_regn_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_final_index_sum_regn_Update/ack
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_base_plus_offset/$entry
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_base_plus_offset/$exit
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_base_plus_offset/sum_rename_req
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2488_base_plus_offset/sum_rename_ack
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_request/$entry
      -- CP-element group 370: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_request/req
      -- 
    ack_4500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2488_index_offset_ack_1, ack => zeropad3D_CP_676_elements(370)); -- 
    req_4509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(370), ack => addr_of_2489_final_reg_req_0); -- 
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_request/$exit
      -- CP-element group 371: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_request/ack
      -- 
    ack_4510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2489_final_reg_ack_0, ack => zeropad3D_CP_676_elements(371)); -- 
    -- CP-element group 372:  join  fork  transition  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	349 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (24) 
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_complete/$exit
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2489_complete/ack
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_sample_start_
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_base_address_calculated
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_word_address_calculated
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_root_address_calculated
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_base_address_resized
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_base_addr_resize/$entry
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_base_addr_resize/$exit
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_base_addr_resize/base_resize_req
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_base_addr_resize/base_resize_ack
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_base_plus_offset/$entry
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_base_plus_offset/$exit
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_base_plus_offset/sum_rename_req
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_base_plus_offset/sum_rename_ack
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_word_addrgen/$entry
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_word_addrgen/$exit
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_word_addrgen/root_register_req
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_word_addrgen/root_register_ack
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Sample/word_access_start/$entry
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Sample/word_access_start/word_0/$entry
      -- CP-element group 372: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Sample/word_access_start/word_0/rr
      -- 
    ack_4515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2489_final_reg_ack_1, ack => zeropad3D_CP_676_elements(372)); -- 
    rr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(372), ack => ptr_deref_2493_load_0_req_0); -- 
    -- CP-element group 373:  transition  input  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373:  members (5) 
      -- CP-element group 373: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_sample_completed_
      -- CP-element group 373: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Sample/$exit
      -- CP-element group 373: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Sample/word_access_start/$exit
      -- CP-element group 373: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Sample/word_access_start/word_0/$exit
      -- CP-element group 373: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Sample/word_access_start/word_0/ra
      -- 
    ra_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2493_load_0_ack_0, ack => zeropad3D_CP_676_elements(373)); -- 
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	349 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	381 
    -- CP-element group 374:  members (9) 
      -- CP-element group 374: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_update_completed_
      -- CP-element group 374: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/$exit
      -- CP-element group 374: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/word_access_complete/$exit
      -- CP-element group 374: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/word_access_complete/word_0/$exit
      -- CP-element group 374: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/word_access_complete/word_0/ca
      -- CP-element group 374: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/ptr_deref_2493_Merge/$entry
      -- CP-element group 374: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/ptr_deref_2493_Merge/$exit
      -- CP-element group 374: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/ptr_deref_2493_Merge/merge_req
      -- CP-element group 374: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2493_Update/ptr_deref_2493_Merge/merge_ack
      -- 
    ca_4560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2493_load_0_ack_1, ack => zeropad3D_CP_676_elements(374)); -- 
    -- CP-element group 375:  transition  input  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	366 
    -- CP-element group 375: successors 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_Sample/ra
      -- 
    ra_4574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2507_inst_ack_0, ack => zeropad3D_CP_676_elements(375)); -- 
    -- CP-element group 376:  transition  input  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	349 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (16) 
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/type_cast_2507_Update/ca
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_resized_1
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_scaled_1
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_computed_1
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_resize_1/$entry
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_resize_1/$exit
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_resize_1/index_resize_req
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_resize_1/index_resize_ack
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_scale_1/$entry
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_scale_1/$exit
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_scale_1/scale_rename_req
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_index_scale_1/scale_rename_ack
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_final_index_sum_regn_Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_final_index_sum_regn_Sample/req
      -- 
    ca_4579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2507_inst_ack_1, ack => zeropad3D_CP_676_elements(376)); -- 
    req_4604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(376), ack => array_obj_ref_2513_index_offset_req_0); -- 
    -- CP-element group 377:  transition  input  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	384 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_final_index_sum_regn_sample_complete
      -- CP-element group 377: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_final_index_sum_regn_Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_final_index_sum_regn_Sample/ack
      -- 
    ack_4605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2513_index_offset_ack_0, ack => zeropad3D_CP_676_elements(377)); -- 
    -- CP-element group 378:  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	349 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (11) 
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_root_address_calculated
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_offset_calculated
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_final_index_sum_regn_Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_final_index_sum_regn_Update/ack
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_base_plus_offset/$entry
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_base_plus_offset/$exit
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_base_plus_offset/sum_rename_req
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/array_obj_ref_2513_base_plus_offset/sum_rename_ack
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_request/$entry
      -- CP-element group 378: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_request/req
      -- 
    ack_4610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2513_index_offset_ack_1, ack => zeropad3D_CP_676_elements(378)); -- 
    req_4619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(378), ack => addr_of_2514_final_reg_req_0); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_sample_completed_
      -- CP-element group 379: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_request/$exit
      -- CP-element group 379: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_request/ack
      -- 
    ack_4620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2514_final_reg_ack_0, ack => zeropad3D_CP_676_elements(379)); -- 
    -- CP-element group 380:  fork  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	349 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (19) 
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_update_completed_
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_complete/$exit
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/addr_of_2514_complete/ack
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_base_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_word_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_root_address_calculated
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_base_address_resized
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_base_addr_resize/$entry
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_base_addr_resize/$exit
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_base_addr_resize/base_resize_req
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_base_addr_resize/base_resize_ack
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_base_plus_offset/$entry
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_base_plus_offset/$exit
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_base_plus_offset/sum_rename_req
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_base_plus_offset/sum_rename_ack
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_word_addrgen/$entry
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_word_addrgen/$exit
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_word_addrgen/root_register_req
      -- CP-element group 380: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_word_addrgen/root_register_ack
      -- 
    ack_4625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2514_final_reg_ack_1, ack => zeropad3D_CP_676_elements(380)); -- 
    -- CP-element group 381:  join  transition  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	374 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (9) 
      -- CP-element group 381: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_sample_start_
      -- CP-element group 381: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/$entry
      -- CP-element group 381: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/ptr_deref_2517_Split/$entry
      -- CP-element group 381: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/ptr_deref_2517_Split/$exit
      -- CP-element group 381: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/ptr_deref_2517_Split/split_req
      -- CP-element group 381: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/ptr_deref_2517_Split/split_ack
      -- CP-element group 381: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/word_access_start/$entry
      -- CP-element group 381: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/word_access_start/word_0/$entry
      -- CP-element group 381: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/word_access_start/word_0/rr
      -- 
    rr_4663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(381), ack => ptr_deref_2517_store_0_req_0); -- 
    zeropad3D_cp_element_group_381: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_381"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(374) & zeropad3D_CP_676_elements(380);
      gj_zeropad3D_cp_element_group_381 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(381), clk => clk, reset => reset); --
    end block;
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382:  members (5) 
      -- CP-element group 382: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/word_access_start/$exit
      -- CP-element group 382: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/word_access_start/word_0/$exit
      -- CP-element group 382: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Sample/word_access_start/word_0/ra
      -- 
    ra_4664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2517_store_0_ack_0, ack => zeropad3D_CP_676_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	349 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (5) 
      -- CP-element group 383: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Update/word_access_complete/$exit
      -- CP-element group 383: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Update/word_access_complete/word_0/$exit
      -- CP-element group 383: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/ptr_deref_2517_Update/word_access_complete/word_0/ca
      -- 
    ca_4675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2517_store_0_ack_1, ack => zeropad3D_CP_676_elements(383)); -- 
    -- CP-element group 384:  join  transition  place  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	369 
    -- CP-element group 384: 	377 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	791 
    -- CP-element group 384:  members (5) 
      -- CP-element group 384: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519__exit__
      -- CP-element group 384: 	 branch_block_stmt_223/ifx_xelse1025_ifx_xend1073
      -- CP-element group 384: 	 branch_block_stmt_223/assign_stmt_2419_to_assign_stmt_2519/$exit
      -- CP-element group 384: 	 branch_block_stmt_223/ifx_xelse1025_ifx_xend1073_PhiReq/$entry
      -- CP-element group 384: 	 branch_block_stmt_223/ifx_xelse1025_ifx_xend1073_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(369) & zeropad3D_CP_676_elements(377) & zeropad3D_CP_676_elements(383);
      gj_zeropad3D_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	791 
    -- CP-element group 385: successors 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_sample_completed_
      -- CP-element group 385: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_Sample/$exit
      -- CP-element group 385: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_Sample/ra
      -- 
    ra_4687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2525_inst_ack_0, ack => zeropad3D_CP_676_elements(385)); -- 
    -- CP-element group 386:  branch  transition  place  input  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	791 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386: 	388 
    -- CP-element group 386:  members (13) 
      -- CP-element group 386: 	 branch_block_stmt_223/if_stmt_2540__entry__
      -- CP-element group 386: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539__exit__
      -- CP-element group 386: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/$exit
      -- CP-element group 386: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_update_completed_
      -- CP-element group 386: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_Update/$exit
      -- CP-element group 386: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_Update/ca
      -- CP-element group 386: 	 branch_block_stmt_223/if_stmt_2540_dead_link/$entry
      -- CP-element group 386: 	 branch_block_stmt_223/if_stmt_2540_eval_test/$entry
      -- CP-element group 386: 	 branch_block_stmt_223/if_stmt_2540_eval_test/$exit
      -- CP-element group 386: 	 branch_block_stmt_223/if_stmt_2540_eval_test/branch_req
      -- CP-element group 386: 	 branch_block_stmt_223/R_cmp1081_2541_place
      -- CP-element group 386: 	 branch_block_stmt_223/if_stmt_2540_if_link/$entry
      -- CP-element group 386: 	 branch_block_stmt_223/if_stmt_2540_else_link/$entry
      -- 
    ca_4692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2525_inst_ack_1, ack => zeropad3D_CP_676_elements(386)); -- 
    branch_req_4700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(386), ack => if_stmt_2540_branch_req_0); -- 
    -- CP-element group 387:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	800 
    -- CP-element group 387: 	801 
    -- CP-element group 387: 	803 
    -- CP-element group 387: 	804 
    -- CP-element group 387: 	806 
    -- CP-element group 387: 	807 
    -- CP-element group 387:  members (40) 
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126
      -- CP-element group 387: 	 branch_block_stmt_223/assign_stmt_2552__exit__
      -- CP-element group 387: 	 branch_block_stmt_223/assign_stmt_2552__entry__
      -- CP-element group 387: 	 branch_block_stmt_223/merge_stmt_2546__exit__
      -- CP-element group 387: 	 branch_block_stmt_223/if_stmt_2540_if_link/$exit
      -- CP-element group 387: 	 branch_block_stmt_223/if_stmt_2540_if_link/if_choice_transition
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xend1073_ifx_xthen1083
      -- CP-element group 387: 	 branch_block_stmt_223/assign_stmt_2552/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/assign_stmt_2552/$exit
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xend1073_ifx_xthen1083_PhiReq/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xend1073_ifx_xthen1083_PhiReq/$exit
      -- CP-element group 387: 	 branch_block_stmt_223/merge_stmt_2546_PhiReqMerge
      -- CP-element group 387: 	 branch_block_stmt_223/merge_stmt_2546_PhiAck/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/merge_stmt_2546_PhiAck/$exit
      -- CP-element group 387: 	 branch_block_stmt_223/merge_stmt_2546_PhiAck/dummy
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Update/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Update/cr
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/SplitProtocol/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/SplitProtocol/Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/SplitProtocol/Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/SplitProtocol/Update/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/SplitProtocol/Update/cr
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/SplitProtocol/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/SplitProtocol/Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/SplitProtocol/Sample/rr
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/SplitProtocol/Update/$entry
      -- CP-element group 387: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2540_branch_ack_1, ack => zeropad3D_CP_676_elements(387)); -- 
    rr_8316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(387), ack => type_cast_2607_inst_req_0); -- 
    cr_8321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(387), ack => type_cast_2607_inst_req_1); -- 
    rr_8339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(387), ack => type_cast_2614_inst_req_0); -- 
    cr_8344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(387), ack => type_cast_2614_inst_req_1); -- 
    rr_8362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(387), ack => type_cast_2620_inst_req_0); -- 
    cr_8367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(387), ack => type_cast_2620_inst_req_1); -- 
    -- CP-element group 388:  fork  transition  place  input  output  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	386 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	389 
    -- CP-element group 388: 	390 
    -- CP-element group 388: 	392 
    -- CP-element group 388: 	394 
    -- CP-element group 388:  members (24) 
      -- CP-element group 388: 	 branch_block_stmt_223/merge_stmt_2554__exit__
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596__entry__
      -- CP-element group 388: 	 branch_block_stmt_223/if_stmt_2540_else_link/$exit
      -- CP-element group 388: 	 branch_block_stmt_223/if_stmt_2540_else_link/else_choice_transition
      -- CP-element group 388: 	 branch_block_stmt_223/ifx_xend1073_ifx_xelse1088
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/$entry
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_sample_start_
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_update_start_
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_Sample/$entry
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_Sample/rr
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_Update/$entry
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_Update/cr
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_update_start_
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_Update/$entry
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_Update/cr
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_update_start_
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_Update/$entry
      -- CP-element group 388: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_Update/cr
      -- CP-element group 388: 	 branch_block_stmt_223/ifx_xend1073_ifx_xelse1088_PhiReq/$entry
      -- CP-element group 388: 	 branch_block_stmt_223/ifx_xend1073_ifx_xelse1088_PhiReq/$exit
      -- CP-element group 388: 	 branch_block_stmt_223/merge_stmt_2554_PhiReqMerge
      -- CP-element group 388: 	 branch_block_stmt_223/merge_stmt_2554_PhiAck/$entry
      -- CP-element group 388: 	 branch_block_stmt_223/merge_stmt_2554_PhiAck/$exit
      -- CP-element group 388: 	 branch_block_stmt_223/merge_stmt_2554_PhiAck/dummy
      -- 
    else_choice_transition_4709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2540_branch_ack_0, ack => zeropad3D_CP_676_elements(388)); -- 
    rr_4725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(388), ack => type_cast_2564_inst_req_0); -- 
    cr_4730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(388), ack => type_cast_2564_inst_req_1); -- 
    cr_4744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(388), ack => type_cast_2573_inst_req_1); -- 
    cr_4758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(388), ack => type_cast_2590_inst_req_1); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	388 
    -- CP-element group 389: successors 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_sample_completed_
      -- CP-element group 389: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_Sample/ra
      -- 
    ra_4726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2564_inst_ack_0, ack => zeropad3D_CP_676_elements(389)); -- 
    -- CP-element group 390:  transition  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	388 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (6) 
      -- CP-element group 390: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_update_completed_
      -- CP-element group 390: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2564_Update/ca
      -- CP-element group 390: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_sample_start_
      -- CP-element group 390: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_Sample/rr
      -- 
    ca_4731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2564_inst_ack_1, ack => zeropad3D_CP_676_elements(390)); -- 
    rr_4739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(390), ack => type_cast_2573_inst_req_0); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_sample_completed_
      -- CP-element group 391: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_Sample/$exit
      -- CP-element group 391: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_Sample/ra
      -- 
    ra_4740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2573_inst_ack_0, ack => zeropad3D_CP_676_elements(391)); -- 
    -- CP-element group 392:  transition  input  output  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	388 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392:  members (6) 
      -- CP-element group 392: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_update_completed_
      -- CP-element group 392: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_Update/$exit
      -- CP-element group 392: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2573_Update/ca
      -- CP-element group 392: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_sample_start_
      -- CP-element group 392: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_Sample/$entry
      -- CP-element group 392: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_Sample/rr
      -- 
    ca_4745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2573_inst_ack_1, ack => zeropad3D_CP_676_elements(392)); -- 
    rr_4753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(392), ack => type_cast_2590_inst_req_0); -- 
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_sample_completed_
      -- CP-element group 393: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_Sample/$exit
      -- CP-element group 393: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_Sample/ra
      -- 
    ra_4754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2590_inst_ack_0, ack => zeropad3D_CP_676_elements(393)); -- 
    -- CP-element group 394:  branch  transition  place  input  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	388 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394: 	396 
    -- CP-element group 394:  members (13) 
      -- CP-element group 394: 	 branch_block_stmt_223/if_stmt_2597__entry__
      -- CP-element group 394: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596__exit__
      -- CP-element group 394: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/$exit
      -- CP-element group 394: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_update_completed_
      -- CP-element group 394: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_Update/$exit
      -- CP-element group 394: 	 branch_block_stmt_223/assign_stmt_2560_to_assign_stmt_2596/type_cast_2590_Update/ca
      -- CP-element group 394: 	 branch_block_stmt_223/if_stmt_2597_dead_link/$entry
      -- CP-element group 394: 	 branch_block_stmt_223/if_stmt_2597_eval_test/$entry
      -- CP-element group 394: 	 branch_block_stmt_223/if_stmt_2597_eval_test/$exit
      -- CP-element group 394: 	 branch_block_stmt_223/if_stmt_2597_eval_test/branch_req
      -- CP-element group 394: 	 branch_block_stmt_223/R_cmp1117_2598_place
      -- CP-element group 394: 	 branch_block_stmt_223/if_stmt_2597_if_link/$entry
      -- CP-element group 394: 	 branch_block_stmt_223/if_stmt_2597_else_link/$entry
      -- 
    ca_4759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2590_inst_ack_1, ack => zeropad3D_CP_676_elements(394)); -- 
    branch_req_4767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(394), ack => if_stmt_2597_branch_req_0); -- 
    -- CP-element group 395:  fork  transition  place  input  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	397 
    -- CP-element group 395: 	398 
    -- CP-element group 395: 	400 
    -- CP-element group 395:  members (27) 
      -- CP-element group 395: 	 branch_block_stmt_223/merge_stmt_2625__exit__
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658__entry__
      -- CP-element group 395: 	 branch_block_stmt_223/if_stmt_2597_if_link/$exit
      -- CP-element group 395: 	 branch_block_stmt_223/if_stmt_2597_if_link/if_choice_transition
      -- CP-element group 395: 	 branch_block_stmt_223/ifx_xelse1088_whilex_xend1127
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/$entry
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_sample_start_
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_update_start_
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_word_address_calculated
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_root_address_calculated
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Sample/$entry
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Sample/word_access_start/$entry
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Sample/word_access_start/word_0/$entry
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Sample/word_access_start/word_0/rr
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/$entry
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/word_access_complete/$entry
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/word_access_complete/word_0/$entry
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/word_access_complete/word_0/cr
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_update_start_
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_Update/$entry
      -- CP-element group 395: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_Update/cr
      -- CP-element group 395: 	 branch_block_stmt_223/ifx_xelse1088_whilex_xend1127_PhiReq/$entry
      -- CP-element group 395: 	 branch_block_stmt_223/ifx_xelse1088_whilex_xend1127_PhiReq/$exit
      -- CP-element group 395: 	 branch_block_stmt_223/merge_stmt_2625_PhiReqMerge
      -- CP-element group 395: 	 branch_block_stmt_223/merge_stmt_2625_PhiAck/$entry
      -- CP-element group 395: 	 branch_block_stmt_223/merge_stmt_2625_PhiAck/$exit
      -- CP-element group 395: 	 branch_block_stmt_223/merge_stmt_2625_PhiAck/dummy
      -- 
    if_choice_transition_4772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2597_branch_ack_1, ack => zeropad3D_CP_676_elements(395)); -- 
    rr_4797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(395), ack => LOAD_pad_2627_load_0_req_0); -- 
    cr_4808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(395), ack => LOAD_pad_2627_load_0_req_1); -- 
    cr_4827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(395), ack => type_cast_2631_inst_req_1); -- 
    -- CP-element group 396:  fork  transition  place  input  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	394 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	792 
    -- CP-element group 396: 	793 
    -- CP-element group 396: 	794 
    -- CP-element group 396: 	796 
    -- CP-element group 396: 	797 
    -- CP-element group 396:  members (22) 
      -- CP-element group 396: 	 branch_block_stmt_223/if_stmt_2597_else_link/$exit
      -- CP-element group 396: 	 branch_block_stmt_223/if_stmt_2597_else_link/else_choice_transition
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2604/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/SplitProtocol/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/SplitProtocol/Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/SplitProtocol/Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/SplitProtocol/Update/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/SplitProtocol/Update/cr
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/SplitProtocol/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/SplitProtocol/Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/SplitProtocol/Sample/rr
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/SplitProtocol/Update/$entry
      -- CP-element group 396: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2597_branch_ack_0, ack => zeropad3D_CP_676_elements(396)); -- 
    rr_8267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(396), ack => type_cast_2616_inst_req_0); -- 
    cr_8272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(396), ack => type_cast_2616_inst_req_1); -- 
    rr_8290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(396), ack => type_cast_2622_inst_req_0); -- 
    cr_8295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(396), ack => type_cast_2622_inst_req_1); -- 
    -- CP-element group 397:  transition  input  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	395 
    -- CP-element group 397: successors 
    -- CP-element group 397:  members (5) 
      -- CP-element group 397: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_sample_completed_
      -- CP-element group 397: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Sample/$exit
      -- CP-element group 397: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Sample/word_access_start/$exit
      -- CP-element group 397: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Sample/word_access_start/word_0/$exit
      -- CP-element group 397: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Sample/word_access_start/word_0/ra
      -- 
    ra_4798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2627_load_0_ack_0, ack => zeropad3D_CP_676_elements(397)); -- 
    -- CP-element group 398:  transition  input  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	395 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (12) 
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_update_completed_
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/$exit
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/word_access_complete/$exit
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/word_access_complete/word_0/$exit
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/word_access_complete/word_0/ca
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/LOAD_pad_2627_Merge/$entry
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/LOAD_pad_2627_Merge/$exit
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/LOAD_pad_2627_Merge/merge_req
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/LOAD_pad_2627_Update/LOAD_pad_2627_Merge/merge_ack
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_Sample/rr
      -- 
    ca_4809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_2627_load_0_ack_1, ack => zeropad3D_CP_676_elements(398)); -- 
    rr_4822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(398), ack => type_cast_2631_inst_req_0); -- 
    -- CP-element group 399:  transition  input  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_sample_completed_
      -- CP-element group 399: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_Sample/$exit
      -- CP-element group 399: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_Sample/ra
      -- 
    ra_4823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2631_inst_ack_0, ack => zeropad3D_CP_676_elements(399)); -- 
    -- CP-element group 400:  fork  transition  place  input  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	395 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	825 
    -- CP-element group 400: 	826 
    -- CP-element group 400: 	827 
    -- CP-element group 400: 	829 
    -- CP-element group 400: 	830 
    -- CP-element group 400:  members (25) 
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191
      -- CP-element group 400: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658__exit__
      -- CP-element group 400: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/$exit
      -- CP-element group 400: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_update_completed_
      -- CP-element group 400: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_Update/$exit
      -- CP-element group 400: 	 branch_block_stmt_223/assign_stmt_2628_to_assign_stmt_2658/type_cast_2631_Update/ca
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2661/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/SplitProtocol/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/SplitProtocol/Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/SplitProtocol/Sample/rr
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/SplitProtocol/Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/SplitProtocol/Update/cr
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/SplitProtocol/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/SplitProtocol/Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/SplitProtocol/Sample/rr
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/SplitProtocol/Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/SplitProtocol/Update/cr
      -- 
    ca_4828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2631_inst_ack_1, ack => zeropad3D_CP_676_elements(400)); -- 
    rr_8483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(400), ack => type_cast_2671_inst_req_0); -- 
    cr_8488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(400), ack => type_cast_2671_inst_req_1); -- 
    rr_8506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(400), ack => type_cast_2677_inst_req_0); -- 
    cr_8511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(400), ack => type_cast_2677_inst_req_1); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	837 
    -- CP-element group 401: successors 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_sample_completed_
      -- CP-element group 401: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_Sample/$exit
      -- CP-element group 401: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_Sample/ra
      -- 
    ra_4840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2684_inst_ack_0, ack => zeropad3D_CP_676_elements(401)); -- 
    -- CP-element group 402:  branch  transition  place  input  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	837 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402: 	404 
    -- CP-element group 402:  members (13) 
      -- CP-element group 402: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710__exit__
      -- CP-element group 402: 	 branch_block_stmt_223/if_stmt_2711__entry__
      -- CP-element group 402: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/$exit
      -- CP-element group 402: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_update_completed_
      -- CP-element group 402: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_Update/$exit
      -- CP-element group 402: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_Update/ca
      -- CP-element group 402: 	 branch_block_stmt_223/if_stmt_2711_dead_link/$entry
      -- CP-element group 402: 	 branch_block_stmt_223/if_stmt_2711_eval_test/$entry
      -- CP-element group 402: 	 branch_block_stmt_223/if_stmt_2711_eval_test/$exit
      -- CP-element group 402: 	 branch_block_stmt_223/if_stmt_2711_eval_test/branch_req
      -- CP-element group 402: 	 branch_block_stmt_223/R_orx_xcond1858_2712_place
      -- CP-element group 402: 	 branch_block_stmt_223/if_stmt_2711_if_link/$entry
      -- CP-element group 402: 	 branch_block_stmt_223/if_stmt_2711_else_link/$entry
      -- 
    ca_4845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2684_inst_ack_1, ack => zeropad3D_CP_676_elements(402)); -- 
    branch_req_4853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(402), ack => if_stmt_2711_branch_req_0); -- 
    -- CP-element group 403:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	405 
    -- CP-element group 403: 	406 
    -- CP-element group 403:  members (18) 
      -- CP-element group 403: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747__entry__
      -- CP-element group 403: 	 branch_block_stmt_223/merge_stmt_2717__exit__
      -- CP-element group 403: 	 branch_block_stmt_223/if_stmt_2711_if_link/$exit
      -- CP-element group 403: 	 branch_block_stmt_223/if_stmt_2711_if_link/if_choice_transition
      -- CP-element group 403: 	 branch_block_stmt_223/whilex_xbody1191_lorx_xlhsx_xfalse1210
      -- CP-element group 403: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/$entry
      -- CP-element group 403: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_update_start_
      -- CP-element group 403: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_Sample/rr
      -- CP-element group 403: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_Update/cr
      -- CP-element group 403: 	 branch_block_stmt_223/merge_stmt_2717_PhiAck/dummy
      -- CP-element group 403: 	 branch_block_stmt_223/merge_stmt_2717_PhiAck/$exit
      -- CP-element group 403: 	 branch_block_stmt_223/whilex_xbody1191_lorx_xlhsx_xfalse1210_PhiReq/$entry
      -- CP-element group 403: 	 branch_block_stmt_223/whilex_xbody1191_lorx_xlhsx_xfalse1210_PhiReq/$exit
      -- CP-element group 403: 	 branch_block_stmt_223/merge_stmt_2717_PhiReqMerge
      -- CP-element group 403: 	 branch_block_stmt_223/merge_stmt_2717_PhiAck/$entry
      -- 
    if_choice_transition_4858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2711_branch_ack_1, ack => zeropad3D_CP_676_elements(403)); -- 
    rr_4875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(403), ack => type_cast_2721_inst_req_0); -- 
    cr_4880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(403), ack => type_cast_2721_inst_req_1); -- 
    -- CP-element group 404:  transition  place  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	402 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	838 
    -- CP-element group 404:  members (5) 
      -- CP-element group 404: 	 branch_block_stmt_223/if_stmt_2711_else_link/$exit
      -- CP-element group 404: 	 branch_block_stmt_223/if_stmt_2711_else_link/else_choice_transition
      -- CP-element group 404: 	 branch_block_stmt_223/whilex_xbody1191_ifx_xthen1227
      -- CP-element group 404: 	 branch_block_stmt_223/whilex_xbody1191_ifx_xthen1227_PhiReq/$entry
      -- CP-element group 404: 	 branch_block_stmt_223/whilex_xbody1191_ifx_xthen1227_PhiReq/$exit
      -- 
    else_choice_transition_4862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2711_branch_ack_0, ack => zeropad3D_CP_676_elements(404)); -- 
    -- CP-element group 405:  transition  input  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	403 
    -- CP-element group 405: successors 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_sample_completed_
      -- CP-element group 405: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_Sample/$exit
      -- CP-element group 405: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_Sample/ra
      -- 
    ra_4876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2721_inst_ack_0, ack => zeropad3D_CP_676_elements(405)); -- 
    -- CP-element group 406:  branch  transition  place  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	403 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406: 	408 
    -- CP-element group 406:  members (13) 
      -- CP-element group 406: 	 branch_block_stmt_223/if_stmt_2748__entry__
      -- CP-element group 406: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747__exit__
      -- CP-element group 406: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/$exit
      -- CP-element group 406: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_update_completed_
      -- CP-element group 406: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_Update/$exit
      -- CP-element group 406: 	 branch_block_stmt_223/assign_stmt_2722_to_assign_stmt_2747/type_cast_2721_Update/ca
      -- CP-element group 406: 	 branch_block_stmt_223/if_stmt_2748_dead_link/$entry
      -- CP-element group 406: 	 branch_block_stmt_223/if_stmt_2748_eval_test/$entry
      -- CP-element group 406: 	 branch_block_stmt_223/if_stmt_2748_eval_test/$exit
      -- CP-element group 406: 	 branch_block_stmt_223/if_stmt_2748_eval_test/branch_req
      -- CP-element group 406: 	 branch_block_stmt_223/R_orx_xcond1859_2749_place
      -- CP-element group 406: 	 branch_block_stmt_223/if_stmt_2748_if_link/$entry
      -- CP-element group 406: 	 branch_block_stmt_223/if_stmt_2748_else_link/$entry
      -- 
    ca_4881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2721_inst_ack_1, ack => zeropad3D_CP_676_elements(406)); -- 
    branch_req_4889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(406), ack => if_stmt_2748_branch_req_0); -- 
    -- CP-element group 407:  fork  transition  place  input  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	423 
    -- CP-element group 407: 	424 
    -- CP-element group 407: 	426 
    -- CP-element group 407: 	428 
    -- CP-element group 407: 	430 
    -- CP-element group 407: 	432 
    -- CP-element group 407: 	434 
    -- CP-element group 407: 	436 
    -- CP-element group 407: 	438 
    -- CP-element group 407: 	441 
    -- CP-element group 407:  members (46) 
      -- CP-element group 407: 	 branch_block_stmt_223/merge_stmt_2812__exit__
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917__entry__
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_update_start_
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_update_start_
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_sample_start_
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_Update/cr
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_update_start_
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_Sample/rr
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_Update/cr
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_Sample/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/if_stmt_2748_if_link/$exit
      -- CP-element group 407: 	 branch_block_stmt_223/if_stmt_2748_if_link/if_choice_transition
      -- CP-element group 407: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1210_ifx_xelse1248
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_final_index_sum_regn_update_start
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_final_index_sum_regn_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_final_index_sum_regn_Update/req
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_complete/req
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_update_start_
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/word_access_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/word_access_complete/word_0/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/word_access_complete/word_0/cr
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_update_start_
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_Update/cr
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_update_start_
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_final_index_sum_regn_update_start
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_final_index_sum_regn_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_final_index_sum_regn_Update/req
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_complete/req
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_update_start_
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Update/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Update/word_access_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Update/word_access_complete/word_0/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Update/word_access_complete/word_0/cr
      -- CP-element group 407: 	 branch_block_stmt_223/merge_stmt_2812_PhiReqMerge
      -- CP-element group 407: 	 branch_block_stmt_223/merge_stmt_2812_PhiAck/dummy
      -- CP-element group 407: 	 branch_block_stmt_223/merge_stmt_2812_PhiAck/$exit
      -- CP-element group 407: 	 branch_block_stmt_223/merge_stmt_2812_PhiAck/$entry
      -- CP-element group 407: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1210_ifx_xelse1248_PhiReq/$exit
      -- CP-element group 407: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1210_ifx_xelse1248_PhiReq/$entry
      -- 
    if_choice_transition_4894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2748_branch_ack_1, ack => zeropad3D_CP_676_elements(407)); -- 
    cr_5057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(407), ack => type_cast_2816_inst_req_1); -- 
    rr_5052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(407), ack => type_cast_2816_inst_req_0); -- 
    cr_5071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(407), ack => type_cast_2880_inst_req_1); -- 
    req_5102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(407), ack => array_obj_ref_2886_index_offset_req_1); -- 
    req_5117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(407), ack => addr_of_2887_final_reg_req_1); -- 
    cr_5162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(407), ack => ptr_deref_2891_load_0_req_1); -- 
    cr_5181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(407), ack => type_cast_2905_inst_req_1); -- 
    req_5212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(407), ack => array_obj_ref_2911_index_offset_req_1); -- 
    req_5227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(407), ack => addr_of_2912_final_reg_req_1); -- 
    cr_5277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(407), ack => ptr_deref_2915_store_0_req_1); -- 
    -- CP-element group 408:  transition  place  input  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	406 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	838 
    -- CP-element group 408:  members (5) 
      -- CP-element group 408: 	 branch_block_stmt_223/if_stmt_2748_else_link/$exit
      -- CP-element group 408: 	 branch_block_stmt_223/if_stmt_2748_else_link/else_choice_transition
      -- CP-element group 408: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1210_ifx_xthen1227
      -- CP-element group 408: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1210_ifx_xthen1227_PhiReq/$entry
      -- CP-element group 408: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1210_ifx_xthen1227_PhiReq/$exit
      -- 
    else_choice_transition_4898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2748_branch_ack_0, ack => zeropad3D_CP_676_elements(408)); -- 
    -- CP-element group 409:  transition  input  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	838 
    -- CP-element group 409: successors 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_sample_completed_
      -- CP-element group 409: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_Sample/$exit
      -- CP-element group 409: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_Sample/ra
      -- 
    ra_4912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2758_inst_ack_0, ack => zeropad3D_CP_676_elements(409)); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	838 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	413 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_update_completed_
      -- CP-element group 410: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_Update/$exit
      -- CP-element group 410: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_Update/ca
      -- 
    ca_4917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2758_inst_ack_1, ack => zeropad3D_CP_676_elements(410)); -- 
    -- CP-element group 411:  transition  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	838 
    -- CP-element group 411: successors 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_Sample/ra
      -- CP-element group 411: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_sample_completed_
      -- CP-element group 411: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_Sample/$exit
      -- 
    ra_4926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2763_inst_ack_0, ack => zeropad3D_CP_676_elements(411)); -- 
    -- CP-element group 412:  transition  input  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	838 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_Update/$exit
      -- CP-element group 412: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_Update/ca
      -- CP-element group 412: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_update_completed_
      -- 
    ca_4931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2763_inst_ack_1, ack => zeropad3D_CP_676_elements(412)); -- 
    -- CP-element group 413:  join  transition  output  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	410 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_sample_start_
      -- CP-element group 413: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_Sample/$entry
      -- CP-element group 413: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_Sample/rr
      -- 
    rr_4939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(413), ack => type_cast_2797_inst_req_0); -- 
    zeropad3D_cp_element_group_413: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_413"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(410) & zeropad3D_CP_676_elements(412);
      gj_zeropad3D_cp_element_group_413 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(413), clk => clk, reset => reset); --
    end block;
    -- CP-element group 414:  transition  input  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_sample_completed_
      -- CP-element group 414: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_Sample/$exit
      -- CP-element group 414: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_Sample/ra
      -- 
    ra_4940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2797_inst_ack_0, ack => zeropad3D_CP_676_elements(414)); -- 
    -- CP-element group 415:  transition  input  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	838 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (16) 
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_scale_1/scale_rename_req
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_scale_1/scale_rename_ack
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_final_index_sum_regn_Sample/$entry
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_final_index_sum_regn_Sample/req
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_update_completed_
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_resized_1
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_scaled_1
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_scale_1/$exit
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_scale_1/$entry
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_resize_1/index_resize_ack
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_resize_1/index_resize_req
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_resize_1/$exit
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_resize_1/$entry
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_index_computed_1
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_Update/ca
      -- CP-element group 415: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_Update/$exit
      -- 
    ca_4945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2797_inst_ack_1, ack => zeropad3D_CP_676_elements(415)); -- 
    req_4970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(415), ack => array_obj_ref_2803_index_offset_req_0); -- 
    -- CP-element group 416:  transition  input  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	422 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_final_index_sum_regn_sample_complete
      -- CP-element group 416: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_final_index_sum_regn_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_final_index_sum_regn_Sample/ack
      -- 
    ack_4971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2803_index_offset_ack_0, ack => zeropad3D_CP_676_elements(416)); -- 
    -- CP-element group 417:  transition  input  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	838 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	418 
    -- CP-element group 417:  members (11) 
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_sample_start_
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_base_plus_offset/sum_rename_ack
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_request/$entry
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_final_index_sum_regn_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_final_index_sum_regn_Update/ack
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_base_plus_offset/$entry
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_request/req
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_base_plus_offset/$exit
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_base_plus_offset/sum_rename_req
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_root_address_calculated
      -- CP-element group 417: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_offset_calculated
      -- 
    ack_4976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2803_index_offset_ack_1, ack => zeropad3D_CP_676_elements(417)); -- 
    req_4985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(417), ack => addr_of_2804_final_reg_req_0); -- 
    -- CP-element group 418:  transition  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	417 
    -- CP-element group 418: successors 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_sample_completed_
      -- CP-element group 418: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_request/$exit
      -- CP-element group 418: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_request/ack
      -- 
    ack_4986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2804_final_reg_ack_0, ack => zeropad3D_CP_676_elements(418)); -- 
    -- CP-element group 419:  join  fork  transition  input  output  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	838 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	420 
    -- CP-element group 419:  members (28) 
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_word_addrgen/$entry
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_complete/ack
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_sample_start_
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_base_address_calculated
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_word_address_calculated
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_root_address_calculated
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_base_address_resized
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_base_addr_resize/$entry
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_base_addr_resize/$exit
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_update_completed_
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_word_addrgen/$exit
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_base_addr_resize/base_resize_req
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_word_addrgen/root_register_req
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_word_addrgen/root_register_ack
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/$entry
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/ptr_deref_2807_Split/$entry
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/ptr_deref_2807_Split/$exit
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/ptr_deref_2807_Split/split_req
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_complete/$exit
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_base_plus_offset/sum_rename_ack
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_base_plus_offset/sum_rename_req
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_base_plus_offset/$exit
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/word_access_start/word_0/rr
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/word_access_start/word_0/$entry
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/word_access_start/$entry
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/ptr_deref_2807_Split/split_ack
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_base_plus_offset/$entry
      -- CP-element group 419: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_base_addr_resize/base_resize_ack
      -- 
    ack_4991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2804_final_reg_ack_1, ack => zeropad3D_CP_676_elements(419)); -- 
    rr_5029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(419), ack => ptr_deref_2807_store_0_req_0); -- 
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	419 
    -- CP-element group 420: successors 
    -- CP-element group 420:  members (5) 
      -- CP-element group 420: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_sample_completed_
      -- CP-element group 420: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/$exit
      -- CP-element group 420: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/word_access_start/word_0/ra
      -- CP-element group 420: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/word_access_start/word_0/$exit
      -- CP-element group 420: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Sample/word_access_start/$exit
      -- 
    ra_5030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2807_store_0_ack_0, ack => zeropad3D_CP_676_elements(420)); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	838 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (5) 
      -- CP-element group 421: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Update/$exit
      -- CP-element group 421: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Update/word_access_complete/$exit
      -- CP-element group 421: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_update_completed_
      -- CP-element group 421: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Update/word_access_complete/word_0/$exit
      -- CP-element group 421: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Update/word_access_complete/word_0/ca
      -- 
    ca_5041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2807_store_0_ack_1, ack => zeropad3D_CP_676_elements(421)); -- 
    -- CP-element group 422:  join  transition  place  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	416 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	839 
    -- CP-element group 422:  members (5) 
      -- CP-element group 422: 	 branch_block_stmt_223/ifx_xthen1227_ifx_xend1296
      -- CP-element group 422: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810__exit__
      -- CP-element group 422: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/$exit
      -- CP-element group 422: 	 branch_block_stmt_223/ifx_xthen1227_ifx_xend1296_PhiReq/$exit
      -- CP-element group 422: 	 branch_block_stmt_223/ifx_xthen1227_ifx_xend1296_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_422: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_422"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(416) & zeropad3D_CP_676_elements(421);
      gj_zeropad3D_cp_element_group_422 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(422), clk => clk, reset => reset); --
    end block;
    -- CP-element group 423:  transition  input  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	407 
    -- CP-element group 423: successors 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_Sample/ra
      -- CP-element group 423: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_sample_completed_
      -- CP-element group 423: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_Sample/$exit
      -- 
    ra_5053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2816_inst_ack_0, ack => zeropad3D_CP_676_elements(423)); -- 
    -- CP-element group 424:  fork  transition  input  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	407 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424: 	433 
    -- CP-element group 424:  members (9) 
      -- CP-element group 424: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_Update/ca
      -- CP-element group 424: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_Sample/rr
      -- CP-element group 424: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_Update/$exit
      -- CP-element group 424: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2816_update_completed_
      -- CP-element group 424: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_Sample/rr
      -- 
    ca_5058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2816_inst_ack_1, ack => zeropad3D_CP_676_elements(424)); -- 
    rr_5066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(424), ack => type_cast_2880_inst_req_0); -- 
    rr_5176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(424), ack => type_cast_2905_inst_req_0); -- 
    -- CP-element group 425:  transition  input  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_sample_completed_
      -- CP-element group 425: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_Sample/$exit
      -- CP-element group 425: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_Sample/ra
      -- 
    ra_5067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2880_inst_ack_0, ack => zeropad3D_CP_676_elements(425)); -- 
    -- CP-element group 426:  transition  input  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	407 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426:  members (16) 
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_resize_1/index_resize_ack
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_resize_1/$exit
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_resize_1/index_resize_req
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_scale_1/$entry
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_resized_1
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_scaled_1
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_scale_1/$exit
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_scale_1/scale_rename_req
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_computed_1
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_update_completed_
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_Update/ca
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2880_Update/$exit
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_resize_1/$entry
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_index_scale_1/scale_rename_ack
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_final_index_sum_regn_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_final_index_sum_regn_Sample/req
      -- 
    ca_5072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2880_inst_ack_1, ack => zeropad3D_CP_676_elements(426)); -- 
    req_5097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(426), ack => array_obj_ref_2886_index_offset_req_0); -- 
    -- CP-element group 427:  transition  input  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	442 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_final_index_sum_regn_sample_complete
      -- CP-element group 427: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_final_index_sum_regn_Sample/$exit
      -- CP-element group 427: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_final_index_sum_regn_Sample/ack
      -- 
    ack_5098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2886_index_offset_ack_0, ack => zeropad3D_CP_676_elements(427)); -- 
    -- CP-element group 428:  transition  input  output  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	407 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428:  members (11) 
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_root_address_calculated
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_offset_calculated
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_sample_start_
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_final_index_sum_regn_Update/$exit
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_final_index_sum_regn_Update/ack
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_base_plus_offset/$entry
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_base_plus_offset/$exit
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_base_plus_offset/sum_rename_req
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2886_base_plus_offset/sum_rename_ack
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_request/$entry
      -- CP-element group 428: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_request/req
      -- 
    ack_5103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2886_index_offset_ack_1, ack => zeropad3D_CP_676_elements(428)); -- 
    req_5112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(428), ack => addr_of_2887_final_reg_req_0); -- 
    -- CP-element group 429:  transition  input  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	428 
    -- CP-element group 429: successors 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_sample_completed_
      -- CP-element group 429: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_request/$exit
      -- CP-element group 429: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_request/ack
      -- 
    ack_5113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2887_final_reg_ack_0, ack => zeropad3D_CP_676_elements(429)); -- 
    -- CP-element group 430:  join  fork  transition  input  output  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	407 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	431 
    -- CP-element group 430:  members (24) 
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_update_completed_
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_complete/$exit
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2887_complete/ack
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_base_address_calculated
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_word_address_calculated
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_root_address_calculated
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_base_address_resized
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_base_addr_resize/$entry
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_base_addr_resize/$exit
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_base_addr_resize/base_resize_req
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_base_addr_resize/base_resize_ack
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_base_plus_offset/$entry
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_base_plus_offset/$exit
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_base_plus_offset/sum_rename_req
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_base_plus_offset/sum_rename_ack
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_word_addrgen/$entry
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_word_addrgen/$exit
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_word_addrgen/root_register_req
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_word_addrgen/root_register_ack
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Sample/word_access_start/$entry
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Sample/word_access_start/word_0/$entry
      -- CP-element group 430: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Sample/word_access_start/word_0/rr
      -- 
    ack_5118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2887_final_reg_ack_1, ack => zeropad3D_CP_676_elements(430)); -- 
    rr_5151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(430), ack => ptr_deref_2891_load_0_req_0); -- 
    -- CP-element group 431:  transition  input  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	430 
    -- CP-element group 431: successors 
    -- CP-element group 431:  members (5) 
      -- CP-element group 431: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_sample_completed_
      -- CP-element group 431: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Sample/$exit
      -- CP-element group 431: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Sample/word_access_start/$exit
      -- CP-element group 431: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Sample/word_access_start/word_0/$exit
      -- CP-element group 431: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Sample/word_access_start/word_0/ra
      -- 
    ra_5152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2891_load_0_ack_0, ack => zeropad3D_CP_676_elements(431)); -- 
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	407 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	439 
    -- CP-element group 432:  members (9) 
      -- CP-element group 432: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_update_completed_
      -- CP-element group 432: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/$exit
      -- CP-element group 432: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/word_access_complete/$exit
      -- CP-element group 432: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/word_access_complete/word_0/$exit
      -- CP-element group 432: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/word_access_complete/word_0/ca
      -- CP-element group 432: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/ptr_deref_2891_Merge/$entry
      -- CP-element group 432: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/ptr_deref_2891_Merge/$exit
      -- CP-element group 432: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/ptr_deref_2891_Merge/merge_req
      -- CP-element group 432: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2891_Update/ptr_deref_2891_Merge/merge_ack
      -- 
    ca_5163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2891_load_0_ack_1, ack => zeropad3D_CP_676_elements(432)); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	424 
    -- CP-element group 433: successors 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_sample_completed_
      -- CP-element group 433: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_Sample/$exit
      -- CP-element group 433: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_Sample/ra
      -- 
    ra_5177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2905_inst_ack_0, ack => zeropad3D_CP_676_elements(433)); -- 
    -- CP-element group 434:  transition  input  output  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	407 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	435 
    -- CP-element group 434:  members (16) 
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_update_completed_
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_Update/$exit
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/type_cast_2905_Update/ca
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_resized_1
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_scaled_1
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_computed_1
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_resize_1/$entry
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_resize_1/$exit
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_resize_1/index_resize_req
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_resize_1/index_resize_ack
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_scale_1/$entry
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_scale_1/$exit
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_scale_1/scale_rename_req
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_index_scale_1/scale_rename_ack
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_final_index_sum_regn_Sample/$entry
      -- CP-element group 434: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_final_index_sum_regn_Sample/req
      -- 
    ca_5182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2905_inst_ack_1, ack => zeropad3D_CP_676_elements(434)); -- 
    req_5207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(434), ack => array_obj_ref_2911_index_offset_req_0); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	434 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	442 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_final_index_sum_regn_sample_complete
      -- CP-element group 435: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_final_index_sum_regn_Sample/$exit
      -- CP-element group 435: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_final_index_sum_regn_Sample/ack
      -- 
    ack_5208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2911_index_offset_ack_0, ack => zeropad3D_CP_676_elements(435)); -- 
    -- CP-element group 436:  transition  input  output  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	407 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	437 
    -- CP-element group 436:  members (11) 
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_request/$entry
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_sample_start_
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_root_address_calculated
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_offset_calculated
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_final_index_sum_regn_Update/$exit
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_final_index_sum_regn_Update/ack
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_base_plus_offset/$entry
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_base_plus_offset/$exit
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_base_plus_offset/sum_rename_req
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/array_obj_ref_2911_base_plus_offset/sum_rename_ack
      -- CP-element group 436: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_request/req
      -- 
    ack_5213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2911_index_offset_ack_1, ack => zeropad3D_CP_676_elements(436)); -- 
    req_5222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(436), ack => addr_of_2912_final_reg_req_0); -- 
    -- CP-element group 437:  transition  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	436 
    -- CP-element group 437: successors 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_sample_completed_
      -- CP-element group 437: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_request/$exit
      -- CP-element group 437: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_request/ack
      -- 
    ack_5223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2912_final_reg_ack_0, ack => zeropad3D_CP_676_elements(437)); -- 
    -- CP-element group 438:  fork  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	407 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	439 
    -- CP-element group 438:  members (19) 
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_update_completed_
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_complete/$exit
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/addr_of_2912_complete/ack
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_base_address_calculated
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_word_address_calculated
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_root_address_calculated
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_base_address_resized
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_base_addr_resize/$entry
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_base_addr_resize/$exit
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_base_addr_resize/base_resize_req
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_base_addr_resize/base_resize_ack
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_base_plus_offset/$entry
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_base_plus_offset/$exit
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_base_plus_offset/sum_rename_req
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_base_plus_offset/sum_rename_ack
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_word_addrgen/$entry
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_word_addrgen/$exit
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_word_addrgen/root_register_req
      -- CP-element group 438: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_word_addrgen/root_register_ack
      -- 
    ack_5228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2912_final_reg_ack_1, ack => zeropad3D_CP_676_elements(438)); -- 
    -- CP-element group 439:  join  transition  output  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	432 
    -- CP-element group 439: 	438 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	440 
    -- CP-element group 439:  members (9) 
      -- CP-element group 439: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_sample_start_
      -- CP-element group 439: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/$entry
      -- CP-element group 439: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/ptr_deref_2915_Split/$entry
      -- CP-element group 439: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/ptr_deref_2915_Split/$exit
      -- CP-element group 439: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/ptr_deref_2915_Split/split_req
      -- CP-element group 439: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/ptr_deref_2915_Split/split_ack
      -- CP-element group 439: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/word_access_start/$entry
      -- CP-element group 439: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/word_access_start/word_0/$entry
      -- CP-element group 439: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/word_access_start/word_0/rr
      -- 
    rr_5266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(439), ack => ptr_deref_2915_store_0_req_0); -- 
    zeropad3D_cp_element_group_439: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_439"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(432) & zeropad3D_CP_676_elements(438);
      gj_zeropad3D_cp_element_group_439 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(439), clk => clk, reset => reset); --
    end block;
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	439 
    -- CP-element group 440: successors 
    -- CP-element group 440:  members (5) 
      -- CP-element group 440: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_sample_completed_
      -- CP-element group 440: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/$exit
      -- CP-element group 440: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/word_access_start/$exit
      -- CP-element group 440: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/word_access_start/word_0/$exit
      -- CP-element group 440: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Sample/word_access_start/word_0/ra
      -- 
    ra_5267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2915_store_0_ack_0, ack => zeropad3D_CP_676_elements(440)); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	407 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	442 
    -- CP-element group 441:  members (5) 
      -- CP-element group 441: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_update_completed_
      -- CP-element group 441: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Update/$exit
      -- CP-element group 441: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Update/word_access_complete/$exit
      -- CP-element group 441: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Update/word_access_complete/word_0/$exit
      -- CP-element group 441: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/ptr_deref_2915_Update/word_access_complete/word_0/ca
      -- 
    ca_5278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2915_store_0_ack_1, ack => zeropad3D_CP_676_elements(441)); -- 
    -- CP-element group 442:  join  transition  place  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	427 
    -- CP-element group 442: 	435 
    -- CP-element group 442: 	441 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	839 
    -- CP-element group 442:  members (5) 
      -- CP-element group 442: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917__exit__
      -- CP-element group 442: 	 branch_block_stmt_223/ifx_xelse1248_ifx_xend1296
      -- CP-element group 442: 	 branch_block_stmt_223/assign_stmt_2817_to_assign_stmt_2917/$exit
      -- CP-element group 442: 	 branch_block_stmt_223/ifx_xelse1248_ifx_xend1296_PhiReq/$exit
      -- CP-element group 442: 	 branch_block_stmt_223/ifx_xelse1248_ifx_xend1296_PhiReq/$entry
      -- 
    zeropad3D_cp_element_group_442: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_442"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(427) & zeropad3D_CP_676_elements(435) & zeropad3D_CP_676_elements(441);
      gj_zeropad3D_cp_element_group_442 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(442), clk => clk, reset => reset); --
    end block;
    -- CP-element group 443:  transition  input  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	839 
    -- CP-element group 443: successors 
    -- CP-element group 443:  members (3) 
      -- CP-element group 443: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_sample_completed_
      -- CP-element group 443: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_Sample/$exit
      -- CP-element group 443: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_Sample/ra
      -- 
    ra_5290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2923_inst_ack_0, ack => zeropad3D_CP_676_elements(443)); -- 
    -- CP-element group 444:  branch  transition  place  input  output  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	839 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	445 
    -- CP-element group 444: 	446 
    -- CP-element group 444:  members (13) 
      -- CP-element group 444: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937__exit__
      -- CP-element group 444: 	 branch_block_stmt_223/if_stmt_2938__entry__
      -- CP-element group 444: 	 branch_block_stmt_223/R_cmp1304_2939_place
      -- CP-element group 444: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/$exit
      -- CP-element group 444: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_update_completed_
      -- CP-element group 444: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_Update/$exit
      -- CP-element group 444: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_Update/ca
      -- CP-element group 444: 	 branch_block_stmt_223/if_stmt_2938_dead_link/$entry
      -- CP-element group 444: 	 branch_block_stmt_223/if_stmt_2938_eval_test/$entry
      -- CP-element group 444: 	 branch_block_stmt_223/if_stmt_2938_eval_test/$exit
      -- CP-element group 444: 	 branch_block_stmt_223/if_stmt_2938_eval_test/branch_req
      -- CP-element group 444: 	 branch_block_stmt_223/if_stmt_2938_if_link/$entry
      -- CP-element group 444: 	 branch_block_stmt_223/if_stmt_2938_else_link/$entry
      -- 
    ca_5295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2923_inst_ack_1, ack => zeropad3D_CP_676_elements(444)); -- 
    branch_req_5303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(444), ack => if_stmt_2938_branch_req_0); -- 
    -- CP-element group 445:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	444 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	848 
    -- CP-element group 445: 	849 
    -- CP-element group 445: 	851 
    -- CP-element group 445: 	852 
    -- CP-element group 445: 	854 
    -- CP-element group 445: 	855 
    -- CP-element group 445:  members (40) 
      -- CP-element group 445: 	 branch_block_stmt_223/merge_stmt_2944__exit__
      -- CP-element group 445: 	 branch_block_stmt_223/assign_stmt_2950__entry__
      -- CP-element group 445: 	 branch_block_stmt_223/assign_stmt_2950__exit__
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xend1296_ifx_xthen1306
      -- CP-element group 445: 	 branch_block_stmt_223/if_stmt_2938_if_link/$exit
      -- CP-element group 445: 	 branch_block_stmt_223/if_stmt_2938_if_link/if_choice_transition
      -- CP-element group 445: 	 branch_block_stmt_223/assign_stmt_2950/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/assign_stmt_2950/$exit
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/SplitProtocol/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/SplitProtocol/Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/SplitProtocol/Sample/rr
      -- CP-element group 445: 	 branch_block_stmt_223/merge_stmt_2944_PhiAck/dummy
      -- CP-element group 445: 	 branch_block_stmt_223/merge_stmt_2944_PhiAck/$exit
      -- CP-element group 445: 	 branch_block_stmt_223/merge_stmt_2944_PhiAck/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/merge_stmt_2944_PhiReqMerge
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xend1296_ifx_xthen1306_PhiReq/$exit
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xend1296_ifx_xthen1306_PhiReq/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/SplitProtocol/Update/cr
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/SplitProtocol/Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/SplitProtocol/Update/cr
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/SplitProtocol/Sample/rr
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/SplitProtocol/Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/SplitProtocol/Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/SplitProtocol/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/SplitProtocol/Update/cr
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/SplitProtocol/Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/SplitProtocol/Sample/rr
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/SplitProtocol/Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/SplitProtocol/$entry
      -- CP-element group 445: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/$entry
      -- 
    if_choice_transition_5308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2938_branch_ack_1, ack => zeropad3D_CP_676_elements(445)); -- 
    rr_8689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(445), ack => type_cast_3011_inst_req_0); -- 
    cr_8671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(445), ack => type_cast_3004_inst_req_1); -- 
    cr_8694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(445), ack => type_cast_3011_inst_req_1); -- 
    rr_8666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(445), ack => type_cast_3004_inst_req_0); -- 
    cr_8717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(445), ack => type_cast_3017_inst_req_1); -- 
    rr_8712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(445), ack => type_cast_3017_inst_req_0); -- 
    -- CP-element group 446:  fork  transition  place  input  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	444 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446: 	448 
    -- CP-element group 446: 	450 
    -- CP-element group 446: 	452 
    -- CP-element group 446:  members (24) 
      -- CP-element group 446: 	 branch_block_stmt_223/merge_stmt_2952__exit__
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993__entry__
      -- CP-element group 446: 	 branch_block_stmt_223/ifx_xend1296_ifx_xelse1311
      -- CP-element group 446: 	 branch_block_stmt_223/if_stmt_2938_else_link/$exit
      -- CP-element group 446: 	 branch_block_stmt_223/if_stmt_2938_else_link/else_choice_transition
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/$entry
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_sample_start_
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_update_start_
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_Sample/$entry
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_Sample/rr
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_Update/cr
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_update_start_
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_Update/cr
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_update_start_
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_Update/cr
      -- CP-element group 446: 	 branch_block_stmt_223/merge_stmt_2952_PhiAck/$entry
      -- CP-element group 446: 	 branch_block_stmt_223/merge_stmt_2952_PhiAck/$exit
      -- CP-element group 446: 	 branch_block_stmt_223/merge_stmt_2952_PhiReqMerge
      -- CP-element group 446: 	 branch_block_stmt_223/ifx_xend1296_ifx_xelse1311_PhiReq/$exit
      -- CP-element group 446: 	 branch_block_stmt_223/ifx_xend1296_ifx_xelse1311_PhiReq/$entry
      -- CP-element group 446: 	 branch_block_stmt_223/merge_stmt_2952_PhiAck/dummy
      -- 
    else_choice_transition_5312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2938_branch_ack_0, ack => zeropad3D_CP_676_elements(446)); -- 
    rr_5328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(446), ack => type_cast_2962_inst_req_0); -- 
    cr_5333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(446), ack => type_cast_2962_inst_req_1); -- 
    cr_5347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(446), ack => type_cast_2971_inst_req_1); -- 
    cr_5361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(446), ack => type_cast_2987_inst_req_1); -- 
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_sample_completed_
      -- CP-element group 447: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_Sample/ra
      -- 
    ra_5329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2962_inst_ack_0, ack => zeropad3D_CP_676_elements(447)); -- 
    -- CP-element group 448:  transition  input  output  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	446 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (6) 
      -- CP-element group 448: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_update_completed_
      -- CP-element group 448: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_Update/$exit
      -- CP-element group 448: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2962_Update/ca
      -- CP-element group 448: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_sample_start_
      -- CP-element group 448: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_Sample/$entry
      -- CP-element group 448: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_Sample/rr
      -- 
    ca_5334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2962_inst_ack_1, ack => zeropad3D_CP_676_elements(448)); -- 
    rr_5342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(448), ack => type_cast_2971_inst_req_0); -- 
    -- CP-element group 449:  transition  input  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_sample_completed_
      -- CP-element group 449: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_Sample/$exit
      -- CP-element group 449: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_Sample/ra
      -- 
    ra_5343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2971_inst_ack_0, ack => zeropad3D_CP_676_elements(449)); -- 
    -- CP-element group 450:  transition  input  output  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	446 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (6) 
      -- CP-element group 450: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_update_completed_
      -- CP-element group 450: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_Update/$exit
      -- CP-element group 450: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2971_Update/ca
      -- CP-element group 450: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_sample_start_
      -- CP-element group 450: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_Sample/$entry
      -- CP-element group 450: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_Sample/rr
      -- 
    ca_5348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2971_inst_ack_1, ack => zeropad3D_CP_676_elements(450)); -- 
    rr_5356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(450), ack => type_cast_2987_inst_req_0); -- 
    -- CP-element group 451:  transition  input  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_sample_completed_
      -- CP-element group 451: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_Sample/$exit
      -- CP-element group 451: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_Sample/ra
      -- 
    ra_5357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2987_inst_ack_0, ack => zeropad3D_CP_676_elements(451)); -- 
    -- CP-element group 452:  branch  transition  place  input  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	446 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452: 	454 
    -- CP-element group 452:  members (13) 
      -- CP-element group 452: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993__exit__
      -- CP-element group 452: 	 branch_block_stmt_223/if_stmt_2994__entry__
      -- CP-element group 452: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/$exit
      -- CP-element group 452: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_update_completed_
      -- CP-element group 452: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_Update/$exit
      -- CP-element group 452: 	 branch_block_stmt_223/assign_stmt_2958_to_assign_stmt_2993/type_cast_2987_Update/ca
      -- CP-element group 452: 	 branch_block_stmt_223/if_stmt_2994_dead_link/$entry
      -- CP-element group 452: 	 branch_block_stmt_223/if_stmt_2994_eval_test/$entry
      -- CP-element group 452: 	 branch_block_stmt_223/if_stmt_2994_eval_test/$exit
      -- CP-element group 452: 	 branch_block_stmt_223/if_stmt_2994_eval_test/branch_req
      -- CP-element group 452: 	 branch_block_stmt_223/R_cmp1339_2995_place
      -- CP-element group 452: 	 branch_block_stmt_223/if_stmt_2994_if_link/$entry
      -- CP-element group 452: 	 branch_block_stmt_223/if_stmt_2994_else_link/$entry
      -- 
    ca_5362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2987_inst_ack_1, ack => zeropad3D_CP_676_elements(452)); -- 
    branch_req_5370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(452), ack => if_stmt_2994_branch_req_0); -- 
    -- CP-element group 453:  fork  transition  place  input  output  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	455 
    -- CP-element group 453: 	456 
    -- CP-element group 453: 	458 
    -- CP-element group 453:  members (27) 
      -- CP-element group 453: 	 branch_block_stmt_223/merge_stmt_3022__exit__
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061__entry__
      -- CP-element group 453: 	 branch_block_stmt_223/if_stmt_2994_if_link/$exit
      -- CP-element group 453: 	 branch_block_stmt_223/if_stmt_2994_if_link/if_choice_transition
      -- CP-element group 453: 	 branch_block_stmt_223/ifx_xelse1311_whilex_xend1349
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/$entry
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_sample_start_
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_update_start_
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_word_address_calculated
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_root_address_calculated
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Sample/$entry
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Sample/word_access_start/$entry
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Sample/word_access_start/word_0/$entry
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Sample/word_access_start/word_0/rr
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/$entry
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/word_access_complete/$entry
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/word_access_complete/word_0/$entry
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/word_access_complete/word_0/cr
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_update_start_
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_Update/$entry
      -- CP-element group 453: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_Update/cr
      -- CP-element group 453: 	 branch_block_stmt_223/merge_stmt_3022_PhiAck/$entry
      -- CP-element group 453: 	 branch_block_stmt_223/merge_stmt_3022_PhiAck/$exit
      -- CP-element group 453: 	 branch_block_stmt_223/merge_stmt_3022_PhiAck/dummy
      -- CP-element group 453: 	 branch_block_stmt_223/merge_stmt_3022_PhiReqMerge
      -- CP-element group 453: 	 branch_block_stmt_223/ifx_xelse1311_whilex_xend1349_PhiReq/$exit
      -- CP-element group 453: 	 branch_block_stmt_223/ifx_xelse1311_whilex_xend1349_PhiReq/$entry
      -- 
    if_choice_transition_5375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2994_branch_ack_1, ack => zeropad3D_CP_676_elements(453)); -- 
    rr_5400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(453), ack => LOAD_pad_3030_load_0_req_0); -- 
    cr_5411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(453), ack => LOAD_pad_3030_load_0_req_1); -- 
    cr_5430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(453), ack => type_cast_3034_inst_req_1); -- 
    -- CP-element group 454:  fork  transition  place  input  output  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	452 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	840 
    -- CP-element group 454: 	841 
    -- CP-element group 454: 	842 
    -- CP-element group 454: 	844 
    -- CP-element group 454: 	845 
    -- CP-element group 454:  members (22) 
      -- CP-element group 454: 	 branch_block_stmt_223/if_stmt_2994_else_link/$exit
      -- CP-element group 454: 	 branch_block_stmt_223/if_stmt_2994_else_link/else_choice_transition
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/SplitProtocol/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/SplitProtocol/Sample/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/SplitProtocol/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/SplitProtocol/Sample/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3001/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/SplitProtocol/Update/cr
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/SplitProtocol/Update/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/SplitProtocol/Update/cr
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/SplitProtocol/Sample/rr
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/SplitProtocol/Update/$entry
      -- CP-element group 454: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/SplitProtocol/Sample/rr
      -- 
    else_choice_transition_5379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2994_branch_ack_0, ack => zeropad3D_CP_676_elements(454)); -- 
    cr_8622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(454), ack => type_cast_3013_inst_req_1); -- 
    cr_8645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(454), ack => type_cast_3019_inst_req_1); -- 
    rr_8617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(454), ack => type_cast_3013_inst_req_0); -- 
    rr_8640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(454), ack => type_cast_3019_inst_req_0); -- 
    -- CP-element group 455:  transition  input  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	453 
    -- CP-element group 455: successors 
    -- CP-element group 455:  members (5) 
      -- CP-element group 455: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_sample_completed_
      -- CP-element group 455: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Sample/$exit
      -- CP-element group 455: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Sample/word_access_start/$exit
      -- CP-element group 455: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Sample/word_access_start/word_0/$exit
      -- CP-element group 455: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Sample/word_access_start/word_0/ra
      -- 
    ra_5401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3030_load_0_ack_0, ack => zeropad3D_CP_676_elements(455)); -- 
    -- CP-element group 456:  transition  input  output  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	453 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (12) 
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_update_completed_
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/$exit
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/word_access_complete/$exit
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/word_access_complete/word_0/$exit
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/word_access_complete/word_0/ca
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/LOAD_pad_3030_Merge/$entry
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/LOAD_pad_3030_Merge/$exit
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/LOAD_pad_3030_Merge/merge_req
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/LOAD_pad_3030_Update/LOAD_pad_3030_Merge/merge_ack
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_sample_start_
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_Sample/$entry
      -- CP-element group 456: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_Sample/rr
      -- 
    ca_5412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3030_load_0_ack_1, ack => zeropad3D_CP_676_elements(456)); -- 
    rr_5425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(456), ack => type_cast_3034_inst_req_0); -- 
    -- CP-element group 457:  transition  input  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_sample_completed_
      -- CP-element group 457: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_Sample/$exit
      -- CP-element group 457: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_Sample/ra
      -- 
    ra_5426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3034_inst_ack_0, ack => zeropad3D_CP_676_elements(457)); -- 
    -- CP-element group 458:  fork  transition  place  input  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	453 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	873 
    -- CP-element group 458: 	874 
    -- CP-element group 458: 	875 
    -- CP-element group 458: 	876 
    -- CP-element group 458:  members (19) 
      -- CP-element group 458: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061__exit__
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410
      -- CP-element group 458: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/$exit
      -- CP-element group 458: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_update_completed_
      -- CP-element group 458: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_Update/$exit
      -- CP-element group 458: 	 branch_block_stmt_223/assign_stmt_3028_to_assign_stmt_3061/type_cast_3034_Update/ca
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3077/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3064/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/SplitProtocol/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/SplitProtocol/Sample/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/SplitProtocol/Sample/rr
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/SplitProtocol/Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/SplitProtocol/Update/cr
      -- 
    ca_5431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3034_inst_ack_1, ack => zeropad3D_CP_676_elements(458)); -- 
    rr_8841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(458), ack => type_cast_3076_inst_req_0); -- 
    cr_8846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(458), ack => type_cast_3076_inst_req_1); -- 
    -- CP-element group 459:  transition  input  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	883 
    -- CP-element group 459: successors 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_sample_completed_
      -- CP-element group 459: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_Sample/$exit
      -- CP-element group 459: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_Sample/ra
      -- 
    ra_5443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3088_inst_ack_0, ack => zeropad3D_CP_676_elements(459)); -- 
    -- CP-element group 460:  branch  transition  place  input  output  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	883 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460: 	462 
    -- CP-element group 460:  members (13) 
      -- CP-element group 460: 	 branch_block_stmt_223/if_stmt_3115__entry__
      -- CP-element group 460: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114__exit__
      -- CP-element group 460: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/$exit
      -- CP-element group 460: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_update_completed_
      -- CP-element group 460: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_Update/$exit
      -- CP-element group 460: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_Update/ca
      -- CP-element group 460: 	 branch_block_stmt_223/if_stmt_3115_dead_link/$entry
      -- CP-element group 460: 	 branch_block_stmt_223/if_stmt_3115_eval_test/$entry
      -- CP-element group 460: 	 branch_block_stmt_223/if_stmt_3115_eval_test/$exit
      -- CP-element group 460: 	 branch_block_stmt_223/if_stmt_3115_eval_test/branch_req
      -- CP-element group 460: 	 branch_block_stmt_223/R_orx_xcond1860_3116_place
      -- CP-element group 460: 	 branch_block_stmt_223/if_stmt_3115_if_link/$entry
      -- CP-element group 460: 	 branch_block_stmt_223/if_stmt_3115_else_link/$entry
      -- 
    ca_5448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3088_inst_ack_1, ack => zeropad3D_CP_676_elements(460)); -- 
    branch_req_5456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(460), ack => if_stmt_3115_branch_req_0); -- 
    -- CP-element group 461:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	463 
    -- CP-element group 461: 	464 
    -- CP-element group 461:  members (18) 
      -- CP-element group 461: 	 branch_block_stmt_223/merge_stmt_3121__exit__
      -- CP-element group 461: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151__entry__
      -- CP-element group 461: 	 branch_block_stmt_223/if_stmt_3115_if_link/$exit
      -- CP-element group 461: 	 branch_block_stmt_223/if_stmt_3115_if_link/if_choice_transition
      -- CP-element group 461: 	 branch_block_stmt_223/whilex_xbody1410_lorx_xlhsx_xfalse1427
      -- CP-element group 461: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/$entry
      -- CP-element group 461: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_sample_start_
      -- CP-element group 461: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_update_start_
      -- CP-element group 461: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_Sample/$entry
      -- CP-element group 461: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_Sample/rr
      -- CP-element group 461: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_Update/cr
      -- CP-element group 461: 	 branch_block_stmt_223/whilex_xbody1410_lorx_xlhsx_xfalse1427_PhiReq/$entry
      -- CP-element group 461: 	 branch_block_stmt_223/whilex_xbody1410_lorx_xlhsx_xfalse1427_PhiReq/$exit
      -- CP-element group 461: 	 branch_block_stmt_223/merge_stmt_3121_PhiReqMerge
      -- CP-element group 461: 	 branch_block_stmt_223/merge_stmt_3121_PhiAck/$entry
      -- CP-element group 461: 	 branch_block_stmt_223/merge_stmt_3121_PhiAck/$exit
      -- CP-element group 461: 	 branch_block_stmt_223/merge_stmt_3121_PhiAck/dummy
      -- 
    if_choice_transition_5461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3115_branch_ack_1, ack => zeropad3D_CP_676_elements(461)); -- 
    rr_5478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(461), ack => type_cast_3125_inst_req_0); -- 
    cr_5483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(461), ack => type_cast_3125_inst_req_1); -- 
    -- CP-element group 462:  transition  place  input  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	460 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	884 
    -- CP-element group 462:  members (5) 
      -- CP-element group 462: 	 branch_block_stmt_223/if_stmt_3115_else_link/$exit
      -- CP-element group 462: 	 branch_block_stmt_223/if_stmt_3115_else_link/else_choice_transition
      -- CP-element group 462: 	 branch_block_stmt_223/whilex_xbody1410_ifx_xthen1445
      -- CP-element group 462: 	 branch_block_stmt_223/whilex_xbody1410_ifx_xthen1445_PhiReq/$entry
      -- CP-element group 462: 	 branch_block_stmt_223/whilex_xbody1410_ifx_xthen1445_PhiReq/$exit
      -- 
    else_choice_transition_5465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3115_branch_ack_0, ack => zeropad3D_CP_676_elements(462)); -- 
    -- CP-element group 463:  transition  input  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	461 
    -- CP-element group 463: successors 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_sample_completed_
      -- CP-element group 463: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_Sample/$exit
      -- CP-element group 463: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_Sample/ra
      -- 
    ra_5479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3125_inst_ack_0, ack => zeropad3D_CP_676_elements(463)); -- 
    -- CP-element group 464:  branch  transition  place  input  output  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	461 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	465 
    -- CP-element group 464: 	466 
    -- CP-element group 464:  members (13) 
      -- CP-element group 464: 	 branch_block_stmt_223/if_stmt_3152__entry__
      -- CP-element group 464: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151__exit__
      -- CP-element group 464: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/$exit
      -- CP-element group 464: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_update_completed_
      -- CP-element group 464: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_Update/$exit
      -- CP-element group 464: 	 branch_block_stmt_223/assign_stmt_3126_to_assign_stmt_3151/type_cast_3125_Update/ca
      -- CP-element group 464: 	 branch_block_stmt_223/if_stmt_3152_dead_link/$entry
      -- CP-element group 464: 	 branch_block_stmt_223/if_stmt_3152_eval_test/$entry
      -- CP-element group 464: 	 branch_block_stmt_223/if_stmt_3152_eval_test/$exit
      -- CP-element group 464: 	 branch_block_stmt_223/if_stmt_3152_eval_test/branch_req
      -- CP-element group 464: 	 branch_block_stmt_223/R_orx_xcond1861_3153_place
      -- CP-element group 464: 	 branch_block_stmt_223/if_stmt_3152_if_link/$entry
      -- CP-element group 464: 	 branch_block_stmt_223/if_stmt_3152_else_link/$entry
      -- 
    ca_5484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3125_inst_ack_1, ack => zeropad3D_CP_676_elements(464)); -- 
    branch_req_5492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(464), ack => if_stmt_3152_branch_req_0); -- 
    -- CP-element group 465:  fork  transition  place  input  output  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	464 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	481 
    -- CP-element group 465: 	482 
    -- CP-element group 465: 	484 
    -- CP-element group 465: 	486 
    -- CP-element group 465: 	488 
    -- CP-element group 465: 	490 
    -- CP-element group 465: 	492 
    -- CP-element group 465: 	494 
    -- CP-element group 465: 	496 
    -- CP-element group 465: 	499 
    -- CP-element group 465:  members (46) 
      -- CP-element group 465: 	 branch_block_stmt_223/merge_stmt_3216__exit__
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321__entry__
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_complete/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_complete/req
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_update_start_
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_update_start_
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_Update/cr
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_final_index_sum_regn_Update/req
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Update/word_access_complete/word_0/cr
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Update/word_access_complete/word_0/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Update/word_access_complete/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_final_index_sum_regn_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_update_start_
      -- CP-element group 465: 	 branch_block_stmt_223/if_stmt_3152_if_link/$exit
      -- CP-element group 465: 	 branch_block_stmt_223/if_stmt_3152_if_link/if_choice_transition
      -- CP-element group 465: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1427_ifx_xelse1466
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/word_access_complete/word_0/cr
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/word_access_complete/word_0/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_final_index_sum_regn_update_start
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_update_start_
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_Sample/rr
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_Update/cr
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_update_start_
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_Update/cr
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_update_start_
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_final_index_sum_regn_update_start
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_final_index_sum_regn_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_final_index_sum_regn_Update/req
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_complete/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_complete/req
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_update_start_
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/word_access_complete/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1427_ifx_xelse1466_PhiReq/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1427_ifx_xelse1466_PhiReq/$exit
      -- CP-element group 465: 	 branch_block_stmt_223/merge_stmt_3216_PhiReqMerge
      -- CP-element group 465: 	 branch_block_stmt_223/merge_stmt_3216_PhiAck/$entry
      -- CP-element group 465: 	 branch_block_stmt_223/merge_stmt_3216_PhiAck/$exit
      -- CP-element group 465: 	 branch_block_stmt_223/merge_stmt_3216_PhiAck/dummy
      -- 
    if_choice_transition_5497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3152_branch_ack_1, ack => zeropad3D_CP_676_elements(465)); -- 
    req_5830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(465), ack => addr_of_3316_final_reg_req_1); -- 
    cr_5784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(465), ack => type_cast_3309_inst_req_1); -- 
    req_5815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(465), ack => array_obj_ref_3315_index_offset_req_1); -- 
    cr_5880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(465), ack => ptr_deref_3319_store_0_req_1); -- 
    cr_5765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(465), ack => ptr_deref_3295_load_0_req_1); -- 
    rr_5655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(465), ack => type_cast_3220_inst_req_0); -- 
    cr_5660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(465), ack => type_cast_3220_inst_req_1); -- 
    cr_5674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(465), ack => type_cast_3284_inst_req_1); -- 
    req_5705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(465), ack => array_obj_ref_3290_index_offset_req_1); -- 
    req_5720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(465), ack => addr_of_3291_final_reg_req_1); -- 
    -- CP-element group 466:  transition  place  input  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	464 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	884 
    -- CP-element group 466:  members (5) 
      -- CP-element group 466: 	 branch_block_stmt_223/if_stmt_3152_else_link/$exit
      -- CP-element group 466: 	 branch_block_stmt_223/if_stmt_3152_else_link/else_choice_transition
      -- CP-element group 466: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1427_ifx_xthen1445
      -- CP-element group 466: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1427_ifx_xthen1445_PhiReq/$entry
      -- CP-element group 466: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1427_ifx_xthen1445_PhiReq/$exit
      -- 
    else_choice_transition_5501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3152_branch_ack_0, ack => zeropad3D_CP_676_elements(466)); -- 
    -- CP-element group 467:  transition  input  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	884 
    -- CP-element group 467: successors 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_sample_completed_
      -- CP-element group 467: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_Sample/$exit
      -- CP-element group 467: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_Sample/ra
      -- 
    ra_5515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3162_inst_ack_0, ack => zeropad3D_CP_676_elements(467)); -- 
    -- CP-element group 468:  transition  input  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	884 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	471 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_update_completed_
      -- CP-element group 468: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_Update/$exit
      -- CP-element group 468: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_Update/ca
      -- 
    ca_5520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3162_inst_ack_1, ack => zeropad3D_CP_676_elements(468)); -- 
    -- CP-element group 469:  transition  input  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	884 
    -- CP-element group 469: successors 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_sample_completed_
      -- CP-element group 469: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_Sample/$exit
      -- CP-element group 469: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_Sample/ra
      -- 
    ra_5529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3167_inst_ack_0, ack => zeropad3D_CP_676_elements(469)); -- 
    -- CP-element group 470:  transition  input  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	884 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	471 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_update_completed_
      -- CP-element group 470: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_Update/$exit
      -- CP-element group 470: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_Update/ca
      -- 
    ca_5534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3167_inst_ack_1, ack => zeropad3D_CP_676_elements(470)); -- 
    -- CP-element group 471:  join  transition  output  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	468 
    -- CP-element group 471: 	470 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	472 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_sample_start_
      -- CP-element group 471: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_Sample/$entry
      -- CP-element group 471: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_Sample/rr
      -- 
    rr_5542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(471), ack => type_cast_3201_inst_req_0); -- 
    zeropad3D_cp_element_group_471: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_471"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(468) & zeropad3D_CP_676_elements(470);
      gj_zeropad3D_cp_element_group_471 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(471), clk => clk, reset => reset); --
    end block;
    -- CP-element group 472:  transition  input  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	471 
    -- CP-element group 472: successors 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_sample_completed_
      -- CP-element group 472: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_Sample/$exit
      -- CP-element group 472: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_Sample/ra
      -- 
    ra_5543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3201_inst_ack_0, ack => zeropad3D_CP_676_elements(472)); -- 
    -- CP-element group 473:  transition  input  output  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	884 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473:  members (16) 
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_update_completed_
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_Update/$exit
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_Update/ca
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_resized_1
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_scaled_1
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_computed_1
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_resize_1/$entry
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_resize_1/$exit
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_resize_1/index_resize_req
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_resize_1/index_resize_ack
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_scale_1/$entry
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_scale_1/$exit
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_scale_1/scale_rename_req
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_index_scale_1/scale_rename_ack
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_final_index_sum_regn_Sample/$entry
      -- CP-element group 473: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_final_index_sum_regn_Sample/req
      -- 
    ca_5548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3201_inst_ack_1, ack => zeropad3D_CP_676_elements(473)); -- 
    req_5573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(473), ack => array_obj_ref_3207_index_offset_req_0); -- 
    -- CP-element group 474:  transition  input  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	480 
    -- CP-element group 474:  members (3) 
      -- CP-element group 474: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_final_index_sum_regn_sample_complete
      -- CP-element group 474: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_final_index_sum_regn_Sample/$exit
      -- CP-element group 474: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_final_index_sum_regn_Sample/ack
      -- 
    ack_5574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 474_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3207_index_offset_ack_0, ack => zeropad3D_CP_676_elements(474)); -- 
    -- CP-element group 475:  transition  input  output  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	884 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	476 
    -- CP-element group 475:  members (11) 
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_sample_start_
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_root_address_calculated
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_offset_calculated
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_final_index_sum_regn_Update/$exit
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_final_index_sum_regn_Update/ack
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_base_plus_offset/$entry
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_base_plus_offset/$exit
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_base_plus_offset/sum_rename_req
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_base_plus_offset/sum_rename_ack
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_request/$entry
      -- CP-element group 475: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_request/req
      -- 
    ack_5579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3207_index_offset_ack_1, ack => zeropad3D_CP_676_elements(475)); -- 
    req_5588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(475), ack => addr_of_3208_final_reg_req_0); -- 
    -- CP-element group 476:  transition  input  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	475 
    -- CP-element group 476: successors 
    -- CP-element group 476:  members (3) 
      -- CP-element group 476: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_sample_completed_
      -- CP-element group 476: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_request/$exit
      -- CP-element group 476: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_request/ack
      -- 
    ack_5589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3208_final_reg_ack_0, ack => zeropad3D_CP_676_elements(476)); -- 
    -- CP-element group 477:  join  fork  transition  input  output  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	884 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	478 
    -- CP-element group 477:  members (28) 
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_update_completed_
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_complete/$exit
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_complete/ack
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_sample_start_
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_base_address_calculated
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_word_address_calculated
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_root_address_calculated
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_base_address_resized
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_base_addr_resize/$entry
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_base_addr_resize/$exit
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_base_addr_resize/base_resize_req
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_base_addr_resize/base_resize_ack
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_base_plus_offset/$entry
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_base_plus_offset/$exit
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_base_plus_offset/sum_rename_req
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_base_plus_offset/sum_rename_ack
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_word_addrgen/$entry
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_word_addrgen/$exit
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_word_addrgen/root_register_req
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_word_addrgen/root_register_ack
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/$entry
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/ptr_deref_3211_Split/$entry
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/ptr_deref_3211_Split/$exit
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/ptr_deref_3211_Split/split_req
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/ptr_deref_3211_Split/split_ack
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/word_access_start/$entry
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/word_access_start/word_0/$entry
      -- CP-element group 477: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/word_access_start/word_0/rr
      -- 
    ack_5594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3208_final_reg_ack_1, ack => zeropad3D_CP_676_elements(477)); -- 
    rr_5632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(477), ack => ptr_deref_3211_store_0_req_0); -- 
    -- CP-element group 478:  transition  input  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	477 
    -- CP-element group 478: successors 
    -- CP-element group 478:  members (5) 
      -- CP-element group 478: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_sample_completed_
      -- CP-element group 478: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/$exit
      -- CP-element group 478: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/word_access_start/$exit
      -- CP-element group 478: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/word_access_start/word_0/$exit
      -- CP-element group 478: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Sample/word_access_start/word_0/ra
      -- 
    ra_5633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3211_store_0_ack_0, ack => zeropad3D_CP_676_elements(478)); -- 
    -- CP-element group 479:  transition  input  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	884 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	480 
    -- CP-element group 479:  members (5) 
      -- CP-element group 479: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_update_completed_
      -- CP-element group 479: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Update/$exit
      -- CP-element group 479: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Update/word_access_complete/$exit
      -- CP-element group 479: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Update/word_access_complete/word_0/$exit
      -- CP-element group 479: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Update/word_access_complete/word_0/ca
      -- 
    ca_5644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3211_store_0_ack_1, ack => zeropad3D_CP_676_elements(479)); -- 
    -- CP-element group 480:  join  transition  place  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	474 
    -- CP-element group 480: 	479 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	885 
    -- CP-element group 480:  members (5) 
      -- CP-element group 480: 	 branch_block_stmt_223/ifx_xthen1445_ifx_xend1514
      -- CP-element group 480: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214__exit__
      -- CP-element group 480: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/$exit
      -- CP-element group 480: 	 branch_block_stmt_223/ifx_xthen1445_ifx_xend1514_PhiReq/$entry
      -- CP-element group 480: 	 branch_block_stmt_223/ifx_xthen1445_ifx_xend1514_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_480: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_480"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(474) & zeropad3D_CP_676_elements(479);
      gj_zeropad3D_cp_element_group_480 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(480), clk => clk, reset => reset); --
    end block;
    -- CP-element group 481:  transition  input  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	465 
    -- CP-element group 481: successors 
    -- CP-element group 481:  members (3) 
      -- CP-element group 481: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_sample_completed_
      -- CP-element group 481: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_Sample/$exit
      -- CP-element group 481: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_Sample/ra
      -- 
    ra_5656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3220_inst_ack_0, ack => zeropad3D_CP_676_elements(481)); -- 
    -- CP-element group 482:  fork  transition  input  output  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	465 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	483 
    -- CP-element group 482: 	491 
    -- CP-element group 482:  members (9) 
      -- CP-element group 482: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_update_completed_
      -- CP-element group 482: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_Update/$exit
      -- CP-element group 482: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3220_Update/ca
      -- CP-element group 482: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_Sample/rr
      -- 
    ca_5661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3220_inst_ack_1, ack => zeropad3D_CP_676_elements(482)); -- 
    rr_5669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(482), ack => type_cast_3284_inst_req_0); -- 
    rr_5779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(482), ack => type_cast_3309_inst_req_0); -- 
    -- CP-element group 483:  transition  input  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	482 
    -- CP-element group 483: successors 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_sample_completed_
      -- CP-element group 483: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_Sample/$exit
      -- CP-element group 483: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_Sample/ra
      -- 
    ra_5670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 483_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3284_inst_ack_0, ack => zeropad3D_CP_676_elements(483)); -- 
    -- CP-element group 484:  transition  input  output  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	465 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	485 
    -- CP-element group 484:  members (16) 
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_update_completed_
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_Update/$exit
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3284_Update/ca
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_resized_1
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_scaled_1
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_computed_1
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_resize_1/$entry
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_resize_1/$exit
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_resize_1/index_resize_req
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_resize_1/index_resize_ack
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_scale_1/$entry
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_scale_1/$exit
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_scale_1/scale_rename_req
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_index_scale_1/scale_rename_ack
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_final_index_sum_regn_Sample/$entry
      -- CP-element group 484: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_final_index_sum_regn_Sample/req
      -- 
    ca_5675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3284_inst_ack_1, ack => zeropad3D_CP_676_elements(484)); -- 
    req_5700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(484), ack => array_obj_ref_3290_index_offset_req_0); -- 
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	484 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	500 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_final_index_sum_regn_sample_complete
      -- CP-element group 485: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_final_index_sum_regn_Sample/$exit
      -- CP-element group 485: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_final_index_sum_regn_Sample/ack
      -- 
    ack_5701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3290_index_offset_ack_0, ack => zeropad3D_CP_676_elements(485)); -- 
    -- CP-element group 486:  transition  input  output  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	465 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (11) 
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_sample_start_
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_root_address_calculated
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_offset_calculated
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_final_index_sum_regn_Update/$exit
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_final_index_sum_regn_Update/ack
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_base_plus_offset/$entry
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_base_plus_offset/$exit
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_base_plus_offset/sum_rename_req
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3290_base_plus_offset/sum_rename_ack
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_request/$entry
      -- CP-element group 486: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_request/req
      -- 
    ack_5706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 486_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3290_index_offset_ack_1, ack => zeropad3D_CP_676_elements(486)); -- 
    req_5715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(486), ack => addr_of_3291_final_reg_req_0); -- 
    -- CP-element group 487:  transition  input  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_sample_completed_
      -- CP-element group 487: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_request/$exit
      -- CP-element group 487: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_request/ack
      -- 
    ack_5716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3291_final_reg_ack_0, ack => zeropad3D_CP_676_elements(487)); -- 
    -- CP-element group 488:  join  fork  transition  input  output  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	465 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	489 
    -- CP-element group 488:  members (24) 
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_update_completed_
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_complete/$exit
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3291_complete/ack
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_sample_start_
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_base_address_calculated
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_word_address_calculated
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_root_address_calculated
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_base_address_resized
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_base_addr_resize/$entry
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_base_addr_resize/$exit
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_base_addr_resize/base_resize_req
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_base_addr_resize/base_resize_ack
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_base_plus_offset/$entry
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_base_plus_offset/$exit
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_base_plus_offset/sum_rename_req
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_base_plus_offset/sum_rename_ack
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_word_addrgen/$entry
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_word_addrgen/$exit
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_word_addrgen/root_register_req
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_word_addrgen/root_register_ack
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Sample/$entry
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Sample/word_access_start/$entry
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Sample/word_access_start/word_0/$entry
      -- CP-element group 488: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Sample/word_access_start/word_0/rr
      -- 
    ack_5721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3291_final_reg_ack_1, ack => zeropad3D_CP_676_elements(488)); -- 
    rr_5754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(488), ack => ptr_deref_3295_load_0_req_0); -- 
    -- CP-element group 489:  transition  input  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	488 
    -- CP-element group 489: successors 
    -- CP-element group 489:  members (5) 
      -- CP-element group 489: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_sample_completed_
      -- CP-element group 489: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Sample/$exit
      -- CP-element group 489: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Sample/word_access_start/$exit
      -- CP-element group 489: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Sample/word_access_start/word_0/$exit
      -- CP-element group 489: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Sample/word_access_start/word_0/ra
      -- 
    ra_5755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3295_load_0_ack_0, ack => zeropad3D_CP_676_elements(489)); -- 
    -- CP-element group 490:  transition  input  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	465 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	497 
    -- CP-element group 490:  members (9) 
      -- CP-element group 490: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/ptr_deref_3295_Merge/merge_ack
      -- CP-element group 490: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/ptr_deref_3295_Merge/merge_req
      -- CP-element group 490: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/ptr_deref_3295_Merge/$exit
      -- CP-element group 490: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/ptr_deref_3295_Merge/$entry
      -- CP-element group 490: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/word_access_complete/word_0/ca
      -- CP-element group 490: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/word_access_complete/word_0/$exit
      -- CP-element group 490: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_update_completed_
      -- CP-element group 490: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/$exit
      -- CP-element group 490: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3295_Update/word_access_complete/$exit
      -- 
    ca_5766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 490_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3295_load_0_ack_1, ack => zeropad3D_CP_676_elements(490)); -- 
    -- CP-element group 491:  transition  input  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	482 
    -- CP-element group 491: successors 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_sample_completed_
      -- CP-element group 491: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_Sample/$exit
      -- CP-element group 491: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_Sample/ra
      -- 
    ra_5780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3309_inst_ack_0, ack => zeropad3D_CP_676_elements(491)); -- 
    -- CP-element group 492:  transition  input  output  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	465 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492:  members (16) 
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_resize_1/index_resize_ack
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_scale_1/$entry
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_scale_1/$exit
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_scale_1/scale_rename_req
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_update_completed_
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_scale_1/scale_rename_ack
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_Update/$exit
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_resize_1/index_resize_req
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_resize_1/$exit
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_resize_1/$entry
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_computed_1
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_scaled_1
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_index_resized_1
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/type_cast_3309_Update/ca
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_final_index_sum_regn_Sample/req
      -- CP-element group 492: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_final_index_sum_regn_Sample/$entry
      -- 
    ca_5785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3309_inst_ack_1, ack => zeropad3D_CP_676_elements(492)); -- 
    req_5810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(492), ack => array_obj_ref_3315_index_offset_req_0); -- 
    -- CP-element group 493:  transition  input  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	492 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	500 
    -- CP-element group 493:  members (3) 
      -- CP-element group 493: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_final_index_sum_regn_sample_complete
      -- CP-element group 493: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_final_index_sum_regn_Sample/ack
      -- CP-element group 493: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_final_index_sum_regn_Sample/$exit
      -- 
    ack_5811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3315_index_offset_ack_0, ack => zeropad3D_CP_676_elements(493)); -- 
    -- CP-element group 494:  transition  input  output  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	465 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (11) 
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_final_index_sum_regn_Update/ack
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_base_plus_offset/$entry
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_base_plus_offset/$exit
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_base_plus_offset/sum_rename_req
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_base_plus_offset/sum_rename_ack
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_request/$entry
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_request/req
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_offset_calculated
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_final_index_sum_regn_Update/$exit
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/array_obj_ref_3315_root_address_calculated
      -- CP-element group 494: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_sample_start_
      -- 
    ack_5816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3315_index_offset_ack_1, ack => zeropad3D_CP_676_elements(494)); -- 
    req_5825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(494), ack => addr_of_3316_final_reg_req_0); -- 
    -- CP-element group 495:  transition  input  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_request/$exit
      -- CP-element group 495: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_request/ack
      -- CP-element group 495: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_sample_completed_
      -- 
    ack_5826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3316_final_reg_ack_0, ack => zeropad3D_CP_676_elements(495)); -- 
    -- CP-element group 496:  fork  transition  input  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	465 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	497 
    -- CP-element group 496:  members (19) 
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_base_address_resized
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_complete/$exit
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_complete/ack
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_base_addr_resize/$entry
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_base_addr_resize/$exit
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_base_addr_resize/base_resize_req
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_base_addr_resize/base_resize_ack
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_base_plus_offset/$entry
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_base_plus_offset/$exit
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_root_address_calculated
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_word_address_calculated
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/addr_of_3316_update_completed_
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_base_address_calculated
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_word_addrgen/root_register_ack
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_word_addrgen/root_register_req
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_word_addrgen/$exit
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_word_addrgen/$entry
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_base_plus_offset/sum_rename_ack
      -- CP-element group 496: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_base_plus_offset/sum_rename_req
      -- 
    ack_5831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3316_final_reg_ack_1, ack => zeropad3D_CP_676_elements(496)); -- 
    -- CP-element group 497:  join  transition  output  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	490 
    -- CP-element group 497: 	496 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	498 
    -- CP-element group 497:  members (9) 
      -- CP-element group 497: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_sample_start_
      -- CP-element group 497: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/word_access_start/word_0/rr
      -- CP-element group 497: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/word_access_start/word_0/$entry
      -- CP-element group 497: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/word_access_start/$entry
      -- CP-element group 497: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/ptr_deref_3319_Split/split_ack
      -- CP-element group 497: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/ptr_deref_3319_Split/split_req
      -- CP-element group 497: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/ptr_deref_3319_Split/$exit
      -- CP-element group 497: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/ptr_deref_3319_Split/$entry
      -- CP-element group 497: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/$entry
      -- 
    rr_5869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(497), ack => ptr_deref_3319_store_0_req_0); -- 
    zeropad3D_cp_element_group_497: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_497"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(490) & zeropad3D_CP_676_elements(496);
      gj_zeropad3D_cp_element_group_497 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(497), clk => clk, reset => reset); --
    end block;
    -- CP-element group 498:  transition  input  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	497 
    -- CP-element group 498: successors 
    -- CP-element group 498:  members (5) 
      -- CP-element group 498: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_sample_completed_
      -- CP-element group 498: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/word_access_start/word_0/ra
      -- CP-element group 498: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/word_access_start/word_0/$exit
      -- CP-element group 498: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/word_access_start/$exit
      -- CP-element group 498: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Sample/$exit
      -- 
    ra_5870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3319_store_0_ack_0, ack => zeropad3D_CP_676_elements(498)); -- 
    -- CP-element group 499:  transition  input  bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	465 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	500 
    -- CP-element group 499:  members (5) 
      -- CP-element group 499: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_update_completed_
      -- CP-element group 499: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Update/word_access_complete/word_0/ca
      -- CP-element group 499: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Update/word_access_complete/word_0/$exit
      -- CP-element group 499: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Update/word_access_complete/$exit
      -- CP-element group 499: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/ptr_deref_3319_Update/$exit
      -- 
    ca_5881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3319_store_0_ack_1, ack => zeropad3D_CP_676_elements(499)); -- 
    -- CP-element group 500:  join  transition  place  bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	485 
    -- CP-element group 500: 	493 
    -- CP-element group 500: 	499 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	885 
    -- CP-element group 500:  members (5) 
      -- CP-element group 500: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321__exit__
      -- CP-element group 500: 	 branch_block_stmt_223/ifx_xelse1466_ifx_xend1514
      -- CP-element group 500: 	 branch_block_stmt_223/assign_stmt_3221_to_assign_stmt_3321/$exit
      -- CP-element group 500: 	 branch_block_stmt_223/ifx_xelse1466_ifx_xend1514_PhiReq/$entry
      -- CP-element group 500: 	 branch_block_stmt_223/ifx_xelse1466_ifx_xend1514_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_500: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_500"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(485) & zeropad3D_CP_676_elements(493) & zeropad3D_CP_676_elements(499);
      gj_zeropad3D_cp_element_group_500 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(500), clk => clk, reset => reset); --
    end block;
    -- CP-element group 501:  transition  input  bypass 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	885 
    -- CP-element group 501: successors 
    -- CP-element group 501:  members (3) 
      -- CP-element group 501: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_sample_completed_
      -- CP-element group 501: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_Sample/$exit
      -- CP-element group 501: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_Sample/ra
      -- 
    ra_5893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3327_inst_ack_0, ack => zeropad3D_CP_676_elements(501)); -- 
    -- CP-element group 502:  branch  transition  place  input  output  bypass 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	885 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	503 
    -- CP-element group 502: 	504 
    -- CP-element group 502:  members (13) 
      -- CP-element group 502: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341__exit__
      -- CP-element group 502: 	 branch_block_stmt_223/if_stmt_3342__entry__
      -- CP-element group 502: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/$exit
      -- CP-element group 502: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_update_completed_
      -- CP-element group 502: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_Update/$exit
      -- CP-element group 502: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_Update/ca
      -- CP-element group 502: 	 branch_block_stmt_223/if_stmt_3342_dead_link/$entry
      -- CP-element group 502: 	 branch_block_stmt_223/if_stmt_3342_eval_test/$entry
      -- CP-element group 502: 	 branch_block_stmt_223/if_stmt_3342_eval_test/$exit
      -- CP-element group 502: 	 branch_block_stmt_223/if_stmt_3342_eval_test/branch_req
      -- CP-element group 502: 	 branch_block_stmt_223/if_stmt_3342_if_link/$entry
      -- CP-element group 502: 	 branch_block_stmt_223/if_stmt_3342_else_link/$entry
      -- CP-element group 502: 	 branch_block_stmt_223/R_cmp1522_3343_place
      -- 
    ca_5898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3327_inst_ack_1, ack => zeropad3D_CP_676_elements(502)); -- 
    branch_req_5906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(502), ack => if_stmt_3342_branch_req_0); -- 
    -- CP-element group 503:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	502 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	894 
    -- CP-element group 503: 	895 
    -- CP-element group 503: 	897 
    -- CP-element group 503: 	898 
    -- CP-element group 503: 	900 
    -- CP-element group 503: 	901 
    -- CP-element group 503:  members (40) 
      -- CP-element group 503: 	 branch_block_stmt_223/merge_stmt_3348__exit__
      -- CP-element group 503: 	 branch_block_stmt_223/assign_stmt_3354__entry__
      -- CP-element group 503: 	 branch_block_stmt_223/assign_stmt_3354__exit__
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565
      -- CP-element group 503: 	 branch_block_stmt_223/assign_stmt_3354/$exit
      -- CP-element group 503: 	 branch_block_stmt_223/assign_stmt_3354/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/if_stmt_3342_if_link/if_choice_transition
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xend1514_ifx_xthen1524
      -- CP-element group 503: 	 branch_block_stmt_223/if_stmt_3342_if_link/$exit
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xend1514_ifx_xthen1524_PhiReq/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xend1514_ifx_xthen1524_PhiReq/$exit
      -- CP-element group 503: 	 branch_block_stmt_223/merge_stmt_3348_PhiReqMerge
      -- CP-element group 503: 	 branch_block_stmt_223/merge_stmt_3348_PhiAck/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/merge_stmt_3348_PhiAck/$exit
      -- CP-element group 503: 	 branch_block_stmt_223/merge_stmt_3348_PhiAck/dummy
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/SplitProtocol/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/SplitProtocol/Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/SplitProtocol/Sample/rr
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/SplitProtocol/Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/SplitProtocol/Update/cr
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/SplitProtocol/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/SplitProtocol/Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/SplitProtocol/Sample/rr
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/SplitProtocol/Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/SplitProtocol/Update/cr
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/SplitProtocol/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/SplitProtocol/Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/SplitProtocol/Sample/rr
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/SplitProtocol/Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 503_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3342_branch_ack_1, ack => zeropad3D_CP_676_elements(503)); -- 
    rr_9001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_3424_inst_req_0); -- 
    cr_9006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_3424_inst_req_1); -- 
    rr_9024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_3412_inst_req_0); -- 
    cr_9029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_3412_inst_req_1); -- 
    rr_9047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_3418_inst_req_0); -- 
    cr_9052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(503), ack => type_cast_3418_inst_req_1); -- 
    -- CP-element group 504:  fork  transition  place  input  output  bypass 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	502 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	505 
    -- CP-element group 504: 	506 
    -- CP-element group 504: 	508 
    -- CP-element group 504: 	510 
    -- CP-element group 504:  members (24) 
      -- CP-element group 504: 	 branch_block_stmt_223/merge_stmt_3356__exit__
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398__entry__
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_Sample/$entry
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_Sample/rr
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_Update/cr
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_update_start_
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_Update/cr
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_sample_start_
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/$entry
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_223/if_stmt_3342_else_link/else_choice_transition
      -- CP-element group 504: 	 branch_block_stmt_223/if_stmt_3342_else_link/$exit
      -- CP-element group 504: 	 branch_block_stmt_223/ifx_xend1514_ifx_xelse1529
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_update_start_
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_Update/cr
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_update_start_
      -- CP-element group 504: 	 branch_block_stmt_223/ifx_xend1514_ifx_xelse1529_PhiReq/$entry
      -- CP-element group 504: 	 branch_block_stmt_223/ifx_xend1514_ifx_xelse1529_PhiReq/$exit
      -- CP-element group 504: 	 branch_block_stmt_223/merge_stmt_3356_PhiReqMerge
      -- CP-element group 504: 	 branch_block_stmt_223/merge_stmt_3356_PhiAck/$entry
      -- CP-element group 504: 	 branch_block_stmt_223/merge_stmt_3356_PhiAck/$exit
      -- CP-element group 504: 	 branch_block_stmt_223/merge_stmt_3356_PhiAck/dummy
      -- 
    else_choice_transition_5915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3342_branch_ack_0, ack => zeropad3D_CP_676_elements(504)); -- 
    rr_5931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(504), ack => type_cast_3366_inst_req_0); -- 
    cr_5936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(504), ack => type_cast_3366_inst_req_1); -- 
    cr_5964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(504), ack => type_cast_3392_inst_req_1); -- 
    cr_5950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(504), ack => type_cast_3375_inst_req_1); -- 
    -- CP-element group 505:  transition  input  bypass 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	504 
    -- CP-element group 505: successors 
    -- CP-element group 505:  members (3) 
      -- CP-element group 505: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_Sample/$exit
      -- CP-element group 505: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_Sample/ra
      -- CP-element group 505: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_sample_completed_
      -- 
    ra_5932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3366_inst_ack_0, ack => zeropad3D_CP_676_elements(505)); -- 
    -- CP-element group 506:  transition  input  output  bypass 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	504 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	507 
    -- CP-element group 506:  members (6) 
      -- CP-element group 506: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_Update/$exit
      -- CP-element group 506: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_Update/ca
      -- CP-element group 506: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_sample_start_
      -- CP-element group 506: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3366_update_completed_
      -- CP-element group 506: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_Sample/rr
      -- CP-element group 506: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_Sample/$entry
      -- 
    ca_5937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 506_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3366_inst_ack_1, ack => zeropad3D_CP_676_elements(506)); -- 
    rr_5945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(506), ack => type_cast_3375_inst_req_0); -- 
    -- CP-element group 507:  transition  input  bypass 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	506 
    -- CP-element group 507: successors 
    -- CP-element group 507:  members (3) 
      -- CP-element group 507: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_Sample/ra
      -- CP-element group 507: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_Sample/$exit
      -- CP-element group 507: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_sample_completed_
      -- 
    ra_5946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 507_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3375_inst_ack_0, ack => zeropad3D_CP_676_elements(507)); -- 
    -- CP-element group 508:  transition  input  output  bypass 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	504 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	509 
    -- CP-element group 508:  members (6) 
      -- CP-element group 508: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_Sample/rr
      -- CP-element group 508: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_Sample/$entry
      -- CP-element group 508: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_sample_start_
      -- CP-element group 508: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_Update/ca
      -- CP-element group 508: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_Update/$exit
      -- CP-element group 508: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3375_update_completed_
      -- 
    ca_5951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 508_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3375_inst_ack_1, ack => zeropad3D_CP_676_elements(508)); -- 
    rr_5959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(508), ack => type_cast_3392_inst_req_0); -- 
    -- CP-element group 509:  transition  input  bypass 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	508 
    -- CP-element group 509: successors 
    -- CP-element group 509:  members (3) 
      -- CP-element group 509: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_Sample/ra
      -- CP-element group 509: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_Sample/$exit
      -- CP-element group 509: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_sample_completed_
      -- 
    ra_5960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 509_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3392_inst_ack_0, ack => zeropad3D_CP_676_elements(509)); -- 
    -- CP-element group 510:  branch  transition  place  input  output  bypass 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	504 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	511 
    -- CP-element group 510: 	512 
    -- CP-element group 510:  members (13) 
      -- CP-element group 510: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398__exit__
      -- CP-element group 510: 	 branch_block_stmt_223/if_stmt_3399__entry__
      -- CP-element group 510: 	 branch_block_stmt_223/if_stmt_3399_else_link/$entry
      -- CP-element group 510: 	 branch_block_stmt_223/if_stmt_3399_if_link/$entry
      -- CP-element group 510: 	 branch_block_stmt_223/if_stmt_3399_eval_test/branch_req
      -- CP-element group 510: 	 branch_block_stmt_223/if_stmt_3399_eval_test/$exit
      -- CP-element group 510: 	 branch_block_stmt_223/if_stmt_3399_eval_test/$entry
      -- CP-element group 510: 	 branch_block_stmt_223/if_stmt_3399_dead_link/$entry
      -- CP-element group 510: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_Update/ca
      -- CP-element group 510: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_Update/$exit
      -- CP-element group 510: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/$exit
      -- CP-element group 510: 	 branch_block_stmt_223/R_cmp1556_3400_place
      -- CP-element group 510: 	 branch_block_stmt_223/assign_stmt_3362_to_assign_stmt_3398/type_cast_3392_update_completed_
      -- 
    ca_5965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3392_inst_ack_1, ack => zeropad3D_CP_676_elements(510)); -- 
    branch_req_5973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(510), ack => if_stmt_3399_branch_req_0); -- 
    -- CP-element group 511:  fork  transition  place  input  output  bypass 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	510 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	513 
    -- CP-element group 511: 	514 
    -- CP-element group 511: 	516 
    -- CP-element group 511:  members (27) 
      -- CP-element group 511: 	 branch_block_stmt_223/merge_stmt_3427__exit__
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472__entry__
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/$entry
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_sample_start_
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_update_start_
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_word_address_calculated
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/$entry
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_root_address_calculated
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Sample/$entry
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Sample/word_access_start/word_0/rr
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/word_access_complete/word_0/$entry
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/word_access_complete/word_0/cr
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Sample/word_access_start/word_0/$entry
      -- CP-element group 511: 	 branch_block_stmt_223/if_stmt_3399_if_link/if_choice_transition
      -- CP-element group 511: 	 branch_block_stmt_223/if_stmt_3399_if_link/$exit
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Sample/word_access_start/$entry
      -- CP-element group 511: 	 branch_block_stmt_223/ifx_xelse1529_whilex_xend1566
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_Update/cr
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_Update/$entry
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/word_access_complete/$entry
      -- CP-element group 511: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_update_start_
      -- CP-element group 511: 	 branch_block_stmt_223/ifx_xelse1529_whilex_xend1566_PhiReq/$entry
      -- CP-element group 511: 	 branch_block_stmt_223/ifx_xelse1529_whilex_xend1566_PhiReq/$exit
      -- CP-element group 511: 	 branch_block_stmt_223/merge_stmt_3427_PhiReqMerge
      -- CP-element group 511: 	 branch_block_stmt_223/merge_stmt_3427_PhiAck/$entry
      -- CP-element group 511: 	 branch_block_stmt_223/merge_stmt_3427_PhiAck/$exit
      -- CP-element group 511: 	 branch_block_stmt_223/merge_stmt_3427_PhiAck/dummy
      -- 
    if_choice_transition_5978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 511_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3399_branch_ack_1, ack => zeropad3D_CP_676_elements(511)); -- 
    rr_6003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(511), ack => LOAD_pad_3441_load_0_req_0); -- 
    cr_6014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(511), ack => LOAD_pad_3441_load_0_req_1); -- 
    cr_6033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(511), ack => type_cast_3445_inst_req_1); -- 
    -- CP-element group 512:  fork  transition  place  input  output  bypass 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	510 
    -- CP-element group 512: successors 
    -- CP-element group 512: 	886 
    -- CP-element group 512: 	887 
    -- CP-element group 512: 	889 
    -- CP-element group 512: 	890 
    -- CP-element group 512: 	891 
    -- CP-element group 512:  members (22) 
      -- CP-element group 512: 	 branch_block_stmt_223/if_stmt_3399_else_link/else_choice_transition
      -- CP-element group 512: 	 branch_block_stmt_223/if_stmt_3399_else_link/$exit
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/SplitProtocol/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/SplitProtocol/Sample/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/SplitProtocol/Sample/rr
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/SplitProtocol/Update/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/SplitProtocol/Update/cr
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3406/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/SplitProtocol/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/SplitProtocol/Sample/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/SplitProtocol/Sample/rr
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/SplitProtocol/Update/$entry
      -- CP-element group 512: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 512_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3399_branch_ack_0, ack => zeropad3D_CP_676_elements(512)); -- 
    rr_8944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(512), ack => type_cast_3422_inst_req_0); -- 
    cr_8949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(512), ack => type_cast_3422_inst_req_1); -- 
    rr_8975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(512), ack => type_cast_3416_inst_req_0); -- 
    cr_8980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(512), ack => type_cast_3416_inst_req_1); -- 
    -- CP-element group 513:  transition  input  bypass 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	511 
    -- CP-element group 513: successors 
    -- CP-element group 513:  members (5) 
      -- CP-element group 513: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_sample_completed_
      -- CP-element group 513: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Sample/$exit
      -- CP-element group 513: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Sample/word_access_start/$exit
      -- CP-element group 513: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Sample/word_access_start/word_0/$exit
      -- CP-element group 513: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Sample/word_access_start/word_0/ra
      -- 
    ra_6004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3441_load_0_ack_0, ack => zeropad3D_CP_676_elements(513)); -- 
    -- CP-element group 514:  transition  input  output  bypass 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	511 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	515 
    -- CP-element group 514:  members (12) 
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_update_completed_
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/$exit
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/word_access_complete/$exit
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/word_access_complete/word_0/$exit
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_Sample/rr
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_Sample/$entry
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_sample_start_
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/LOAD_pad_3441_Merge/merge_ack
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/LOAD_pad_3441_Merge/merge_req
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/LOAD_pad_3441_Merge/$exit
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/LOAD_pad_3441_Merge/$entry
      -- CP-element group 514: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/LOAD_pad_3441_Update/word_access_complete/word_0/ca
      -- 
    ca_6015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_pad_3441_load_0_ack_1, ack => zeropad3D_CP_676_elements(514)); -- 
    rr_6028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(514), ack => type_cast_3445_inst_req_0); -- 
    -- CP-element group 515:  transition  input  bypass 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	514 
    -- CP-element group 515: successors 
    -- CP-element group 515:  members (3) 
      -- CP-element group 515: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_Sample/ra
      -- CP-element group 515: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_Sample/$exit
      -- CP-element group 515: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_sample_completed_
      -- 
    ra_6029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 515_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3445_inst_ack_0, ack => zeropad3D_CP_676_elements(515)); -- 
    -- CP-element group 516:  fork  transition  place  input  output  bypass 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	511 
    -- CP-element group 516: successors 
    -- CP-element group 516: 	919 
    -- CP-element group 516: 	920 
    -- CP-element group 516: 	921 
    -- CP-element group 516: 	923 
    -- CP-element group 516: 	924 
    -- CP-element group 516:  members (25) 
      -- CP-element group 516: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472__exit__
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631
      -- CP-element group 516: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/$exit
      -- CP-element group 516: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_Update/ca
      -- CP-element group 516: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_Update/$exit
      -- CP-element group 516: 	 branch_block_stmt_223/assign_stmt_3433_to_assign_stmt_3472/type_cast_3445_update_completed_
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3475/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/SplitProtocol/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/SplitProtocol/Sample/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/SplitProtocol/Sample/rr
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/SplitProtocol/Update/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/SplitProtocol/Update/cr
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/SplitProtocol/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/SplitProtocol/Sample/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/SplitProtocol/Sample/rr
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/SplitProtocol/Update/$entry
      -- CP-element group 516: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/SplitProtocol/Update/cr
      -- 
    ca_6034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 516_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3445_inst_ack_1, ack => zeropad3D_CP_676_elements(516)); -- 
    rr_9168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(516), ack => type_cast_3485_inst_req_0); -- 
    cr_9173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(516), ack => type_cast_3485_inst_req_1); -- 
    rr_9191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(516), ack => type_cast_3491_inst_req_0); -- 
    cr_9196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(516), ack => type_cast_3491_inst_req_1); -- 
    -- CP-element group 517:  transition  input  bypass 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	931 
    -- CP-element group 517: successors 
    -- CP-element group 517:  members (3) 
      -- CP-element group 517: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_Sample/$exit
      -- CP-element group 517: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_Sample/ra
      -- CP-element group 517: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_sample_completed_
      -- 
    ra_6046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3498_inst_ack_0, ack => zeropad3D_CP_676_elements(517)); -- 
    -- CP-element group 518:  branch  transition  place  input  output  bypass 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	931 
    -- CP-element group 518: successors 
    -- CP-element group 518: 	519 
    -- CP-element group 518: 	520 
    -- CP-element group 518:  members (13) 
      -- CP-element group 518: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524__exit__
      -- CP-element group 518: 	 branch_block_stmt_223/if_stmt_3525__entry__
      -- CP-element group 518: 	 branch_block_stmt_223/if_stmt_3525_else_link/$entry
      -- CP-element group 518: 	 branch_block_stmt_223/if_stmt_3525_eval_test/$entry
      -- CP-element group 518: 	 branch_block_stmt_223/if_stmt_3525_eval_test/$exit
      -- CP-element group 518: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_Update/$exit
      -- CP-element group 518: 	 branch_block_stmt_223/if_stmt_3525_eval_test/branch_req
      -- CP-element group 518: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_Update/ca
      -- CP-element group 518: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_update_completed_
      -- CP-element group 518: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/$exit
      -- CP-element group 518: 	 branch_block_stmt_223/R_orx_xcond1862_3526_place
      -- CP-element group 518: 	 branch_block_stmt_223/if_stmt_3525_if_link/$entry
      -- CP-element group 518: 	 branch_block_stmt_223/if_stmt_3525_dead_link/$entry
      -- 
    ca_6051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 518_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3498_inst_ack_1, ack => zeropad3D_CP_676_elements(518)); -- 
    branch_req_6059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(518), ack => if_stmt_3525_branch_req_0); -- 
    -- CP-element group 519:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	518 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	521 
    -- CP-element group 519: 	522 
    -- CP-element group 519:  members (18) 
      -- CP-element group 519: 	 branch_block_stmt_223/merge_stmt_3531__exit__
      -- CP-element group 519: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561__entry__
      -- CP-element group 519: 	 branch_block_stmt_223/whilex_xbody1631_lorx_xlhsx_xfalse1648
      -- CP-element group 519: 	 branch_block_stmt_223/if_stmt_3525_if_link/if_choice_transition
      -- CP-element group 519: 	 branch_block_stmt_223/if_stmt_3525_if_link/$exit
      -- CP-element group 519: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_Update/cr
      -- CP-element group 519: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_Update/$entry
      -- CP-element group 519: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_Sample/rr
      -- CP-element group 519: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_Sample/$entry
      -- CP-element group 519: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_update_start_
      -- CP-element group 519: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_sample_start_
      -- CP-element group 519: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/$entry
      -- CP-element group 519: 	 branch_block_stmt_223/whilex_xbody1631_lorx_xlhsx_xfalse1648_PhiReq/$entry
      -- CP-element group 519: 	 branch_block_stmt_223/whilex_xbody1631_lorx_xlhsx_xfalse1648_PhiReq/$exit
      -- CP-element group 519: 	 branch_block_stmt_223/merge_stmt_3531_PhiReqMerge
      -- CP-element group 519: 	 branch_block_stmt_223/merge_stmt_3531_PhiAck/$entry
      -- CP-element group 519: 	 branch_block_stmt_223/merge_stmt_3531_PhiAck/$exit
      -- CP-element group 519: 	 branch_block_stmt_223/merge_stmt_3531_PhiAck/dummy
      -- 
    if_choice_transition_6064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 519_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3525_branch_ack_1, ack => zeropad3D_CP_676_elements(519)); -- 
    cr_6086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(519), ack => type_cast_3535_inst_req_1); -- 
    rr_6081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(519), ack => type_cast_3535_inst_req_0); -- 
    -- CP-element group 520:  transition  place  input  bypass 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	518 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	932 
    -- CP-element group 520:  members (5) 
      -- CP-element group 520: 	 branch_block_stmt_223/whilex_xbody1631_ifx_xthen1665
      -- CP-element group 520: 	 branch_block_stmt_223/if_stmt_3525_else_link/$exit
      -- CP-element group 520: 	 branch_block_stmt_223/if_stmt_3525_else_link/else_choice_transition
      -- CP-element group 520: 	 branch_block_stmt_223/whilex_xbody1631_ifx_xthen1665_PhiReq/$entry
      -- CP-element group 520: 	 branch_block_stmt_223/whilex_xbody1631_ifx_xthen1665_PhiReq/$exit
      -- 
    else_choice_transition_6068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 520_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3525_branch_ack_0, ack => zeropad3D_CP_676_elements(520)); -- 
    -- CP-element group 521:  transition  input  bypass 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	519 
    -- CP-element group 521: successors 
    -- CP-element group 521:  members (3) 
      -- CP-element group 521: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_Sample/ra
      -- CP-element group 521: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_Sample/$exit
      -- CP-element group 521: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_sample_completed_
      -- 
    ra_6082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3535_inst_ack_0, ack => zeropad3D_CP_676_elements(521)); -- 
    -- CP-element group 522:  branch  transition  place  input  output  bypass 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	519 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	523 
    -- CP-element group 522: 	524 
    -- CP-element group 522:  members (13) 
      -- CP-element group 522: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561__exit__
      -- CP-element group 522: 	 branch_block_stmt_223/if_stmt_3562__entry__
      -- CP-element group 522: 	 branch_block_stmt_223/R_orx_xcond1863_3563_place
      -- CP-element group 522: 	 branch_block_stmt_223/if_stmt_3562_else_link/$entry
      -- CP-element group 522: 	 branch_block_stmt_223/if_stmt_3562_if_link/$entry
      -- CP-element group 522: 	 branch_block_stmt_223/if_stmt_3562_eval_test/branch_req
      -- CP-element group 522: 	 branch_block_stmt_223/if_stmt_3562_eval_test/$exit
      -- CP-element group 522: 	 branch_block_stmt_223/if_stmt_3562_eval_test/$entry
      -- CP-element group 522: 	 branch_block_stmt_223/if_stmt_3562_dead_link/$entry
      -- CP-element group 522: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_Update/ca
      -- CP-element group 522: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_Update/$exit
      -- CP-element group 522: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/type_cast_3535_update_completed_
      -- CP-element group 522: 	 branch_block_stmt_223/assign_stmt_3536_to_assign_stmt_3561/$exit
      -- 
    ca_6087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 522_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3535_inst_ack_1, ack => zeropad3D_CP_676_elements(522)); -- 
    branch_req_6095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(522), ack => if_stmt_3562_branch_req_0); -- 
    -- CP-element group 523:  fork  transition  place  input  output  bypass 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	522 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	539 
    -- CP-element group 523: 	540 
    -- CP-element group 523: 	542 
    -- CP-element group 523: 	544 
    -- CP-element group 523: 	546 
    -- CP-element group 523: 	548 
    -- CP-element group 523: 	550 
    -- CP-element group 523: 	552 
    -- CP-element group 523: 	554 
    -- CP-element group 523: 	557 
    -- CP-element group 523:  members (46) 
      -- CP-element group 523: 	 branch_block_stmt_223/merge_stmt_3626__exit__
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731__entry__
      -- CP-element group 523: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1648_ifx_xelse1686
      -- CP-element group 523: 	 branch_block_stmt_223/if_stmt_3562_if_link/if_choice_transition
      -- CP-element group 523: 	 branch_block_stmt_223/if_stmt_3562_if_link/$exit
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_sample_start_
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_update_start_
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_Sample/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_Sample/rr
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_Update/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_Update/cr
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_update_start_
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_Update/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_Update/cr
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_update_start_
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_final_index_sum_regn_update_start
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_final_index_sum_regn_Update/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_final_index_sum_regn_Update/req
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_complete/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_complete/req
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_update_start_
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/word_access_complete/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/word_access_complete/word_0/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/word_access_complete/word_0/cr
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_update_start_
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_Update/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_Update/cr
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_update_start_
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_final_index_sum_regn_update_start
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_final_index_sum_regn_Update/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_final_index_sum_regn_Update/req
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_complete/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_complete/req
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_update_start_
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Update/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Update/word_access_complete/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Update/word_access_complete/word_0/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Update/word_access_complete/word_0/cr
      -- CP-element group 523: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1648_ifx_xelse1686_PhiReq/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1648_ifx_xelse1686_PhiReq/$exit
      -- CP-element group 523: 	 branch_block_stmt_223/merge_stmt_3626_PhiReqMerge
      -- CP-element group 523: 	 branch_block_stmt_223/merge_stmt_3626_PhiAck/$entry
      -- CP-element group 523: 	 branch_block_stmt_223/merge_stmt_3626_PhiAck/$exit
      -- CP-element group 523: 	 branch_block_stmt_223/merge_stmt_3626_PhiAck/dummy
      -- 
    if_choice_transition_6100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 523_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3562_branch_ack_1, ack => zeropad3D_CP_676_elements(523)); -- 
    rr_6258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => type_cast_3630_inst_req_0); -- 
    cr_6263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => type_cast_3630_inst_req_1); -- 
    cr_6277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => type_cast_3694_inst_req_1); -- 
    req_6308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => array_obj_ref_3700_index_offset_req_1); -- 
    req_6323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => addr_of_3701_final_reg_req_1); -- 
    cr_6368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => ptr_deref_3705_load_0_req_1); -- 
    cr_6387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => type_cast_3719_inst_req_1); -- 
    req_6418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => array_obj_ref_3725_index_offset_req_1); -- 
    req_6433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => addr_of_3726_final_reg_req_1); -- 
    cr_6483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(523), ack => ptr_deref_3729_store_0_req_1); -- 
    -- CP-element group 524:  transition  place  input  bypass 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	522 
    -- CP-element group 524: successors 
    -- CP-element group 524: 	932 
    -- CP-element group 524:  members (5) 
      -- CP-element group 524: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1648_ifx_xthen1665
      -- CP-element group 524: 	 branch_block_stmt_223/if_stmt_3562_else_link/else_choice_transition
      -- CP-element group 524: 	 branch_block_stmt_223/if_stmt_3562_else_link/$exit
      -- CP-element group 524: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1648_ifx_xthen1665_PhiReq/$entry
      -- CP-element group 524: 	 branch_block_stmt_223/lorx_xlhsx_xfalse1648_ifx_xthen1665_PhiReq/$exit
      -- 
    else_choice_transition_6104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3562_branch_ack_0, ack => zeropad3D_CP_676_elements(524)); -- 
    -- CP-element group 525:  transition  input  bypass 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	932 
    -- CP-element group 525: successors 
    -- CP-element group 525:  members (3) 
      -- CP-element group 525: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_sample_completed_
      -- CP-element group 525: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_Sample/$exit
      -- CP-element group 525: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_Sample/ra
      -- 
    ra_6118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 525_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3572_inst_ack_0, ack => zeropad3D_CP_676_elements(525)); -- 
    -- CP-element group 526:  transition  input  bypass 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	932 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	529 
    -- CP-element group 526:  members (3) 
      -- CP-element group 526: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_update_completed_
      -- CP-element group 526: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_Update/ca
      -- CP-element group 526: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_Update/$exit
      -- 
    ca_6123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 526_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3572_inst_ack_1, ack => zeropad3D_CP_676_elements(526)); -- 
    -- CP-element group 527:  transition  input  bypass 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	932 
    -- CP-element group 527: successors 
    -- CP-element group 527:  members (3) 
      -- CP-element group 527: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_sample_completed_
      -- CP-element group 527: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_Sample/ra
      -- CP-element group 527: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_Sample/$exit
      -- 
    ra_6132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 527_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3577_inst_ack_0, ack => zeropad3D_CP_676_elements(527)); -- 
    -- CP-element group 528:  transition  input  bypass 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	932 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	529 
    -- CP-element group 528:  members (3) 
      -- CP-element group 528: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_update_completed_
      -- CP-element group 528: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_Update/ca
      -- CP-element group 528: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_Update/$exit
      -- 
    ca_6137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 528_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3577_inst_ack_1, ack => zeropad3D_CP_676_elements(528)); -- 
    -- CP-element group 529:  join  transition  output  bypass 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	526 
    -- CP-element group 529: 	528 
    -- CP-element group 529: successors 
    -- CP-element group 529: 	530 
    -- CP-element group 529:  members (3) 
      -- CP-element group 529: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_Sample/rr
      -- CP-element group 529: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_Sample/$entry
      -- CP-element group 529: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_sample_start_
      -- 
    rr_6145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(529), ack => type_cast_3611_inst_req_0); -- 
    zeropad3D_cp_element_group_529: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_529"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(526) & zeropad3D_CP_676_elements(528);
      gj_zeropad3D_cp_element_group_529 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(529), clk => clk, reset => reset); --
    end block;
    -- CP-element group 530:  transition  input  bypass 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	529 
    -- CP-element group 530: successors 
    -- CP-element group 530:  members (3) 
      -- CP-element group 530: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_Sample/ra
      -- CP-element group 530: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_Sample/$exit
      -- CP-element group 530: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_sample_completed_
      -- 
    ra_6146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 530_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3611_inst_ack_0, ack => zeropad3D_CP_676_elements(530)); -- 
    -- CP-element group 531:  transition  input  output  bypass 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	932 
    -- CP-element group 531: successors 
    -- CP-element group 531: 	532 
    -- CP-element group 531:  members (16) 
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_Update/ca
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_Update/$exit
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_update_completed_
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_resized_1
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_scaled_1
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_computed_1
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_resize_1/$entry
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_resize_1/$exit
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_resize_1/index_resize_req
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_resize_1/index_resize_ack
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_scale_1/$entry
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_scale_1/$exit
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_scale_1/scale_rename_req
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_index_scale_1/scale_rename_ack
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_final_index_sum_regn_Sample/$entry
      -- CP-element group 531: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_final_index_sum_regn_Sample/req
      -- 
    ca_6151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 531_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3611_inst_ack_1, ack => zeropad3D_CP_676_elements(531)); -- 
    req_6176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(531), ack => array_obj_ref_3617_index_offset_req_0); -- 
    -- CP-element group 532:  transition  input  bypass 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	531 
    -- CP-element group 532: successors 
    -- CP-element group 532: 	538 
    -- CP-element group 532:  members (3) 
      -- CP-element group 532: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_final_index_sum_regn_sample_complete
      -- CP-element group 532: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_final_index_sum_regn_Sample/$exit
      -- CP-element group 532: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_final_index_sum_regn_Sample/ack
      -- 
    ack_6177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 532_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3617_index_offset_ack_0, ack => zeropad3D_CP_676_elements(532)); -- 
    -- CP-element group 533:  transition  input  output  bypass 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	932 
    -- CP-element group 533: successors 
    -- CP-element group 533: 	534 
    -- CP-element group 533:  members (11) 
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_sample_start_
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_root_address_calculated
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_offset_calculated
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_final_index_sum_regn_Update/$exit
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_final_index_sum_regn_Update/ack
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_base_plus_offset/$entry
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_base_plus_offset/$exit
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_base_plus_offset/sum_rename_req
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_base_plus_offset/sum_rename_ack
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_request/$entry
      -- CP-element group 533: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_request/req
      -- 
    ack_6182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 533_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3617_index_offset_ack_1, ack => zeropad3D_CP_676_elements(533)); -- 
    req_6191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(533), ack => addr_of_3618_final_reg_req_0); -- 
    -- CP-element group 534:  transition  input  bypass 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	533 
    -- CP-element group 534: successors 
    -- CP-element group 534:  members (3) 
      -- CP-element group 534: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_sample_completed_
      -- CP-element group 534: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_request/$exit
      -- CP-element group 534: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_request/ack
      -- 
    ack_6192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 534_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3618_final_reg_ack_0, ack => zeropad3D_CP_676_elements(534)); -- 
    -- CP-element group 535:  join  fork  transition  input  output  bypass 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	932 
    -- CP-element group 535: successors 
    -- CP-element group 535: 	536 
    -- CP-element group 535:  members (28) 
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_update_completed_
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_complete/$exit
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_complete/ack
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_sample_start_
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_base_address_calculated
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_word_address_calculated
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_root_address_calculated
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_base_address_resized
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_base_addr_resize/$entry
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_base_addr_resize/$exit
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_base_addr_resize/base_resize_req
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_base_addr_resize/base_resize_ack
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_base_plus_offset/$entry
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_base_plus_offset/$exit
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_base_plus_offset/sum_rename_req
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_base_plus_offset/sum_rename_ack
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_word_addrgen/$entry
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_word_addrgen/$exit
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_word_addrgen/root_register_req
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_word_addrgen/root_register_ack
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/$entry
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/ptr_deref_3621_Split/$entry
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/ptr_deref_3621_Split/$exit
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/ptr_deref_3621_Split/split_req
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/ptr_deref_3621_Split/split_ack
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/word_access_start/$entry
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/word_access_start/word_0/$entry
      -- CP-element group 535: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/word_access_start/word_0/rr
      -- 
    ack_6197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 535_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3618_final_reg_ack_1, ack => zeropad3D_CP_676_elements(535)); -- 
    rr_6235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(535), ack => ptr_deref_3621_store_0_req_0); -- 
    -- CP-element group 536:  transition  input  bypass 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	535 
    -- CP-element group 536: successors 
    -- CP-element group 536:  members (5) 
      -- CP-element group 536: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_sample_completed_
      -- CP-element group 536: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/$exit
      -- CP-element group 536: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/word_access_start/$exit
      -- CP-element group 536: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/word_access_start/word_0/$exit
      -- CP-element group 536: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Sample/word_access_start/word_0/ra
      -- 
    ra_6236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 536_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3621_store_0_ack_0, ack => zeropad3D_CP_676_elements(536)); -- 
    -- CP-element group 537:  transition  input  bypass 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	932 
    -- CP-element group 537: successors 
    -- CP-element group 537: 	538 
    -- CP-element group 537:  members (5) 
      -- CP-element group 537: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_update_completed_
      -- CP-element group 537: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Update/$exit
      -- CP-element group 537: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Update/word_access_complete/$exit
      -- CP-element group 537: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Update/word_access_complete/word_0/$exit
      -- CP-element group 537: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Update/word_access_complete/word_0/ca
      -- 
    ca_6247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 537_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3621_store_0_ack_1, ack => zeropad3D_CP_676_elements(537)); -- 
    -- CP-element group 538:  join  transition  place  bypass 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: 	532 
    -- CP-element group 538: 	537 
    -- CP-element group 538: successors 
    -- CP-element group 538: 	933 
    -- CP-element group 538:  members (5) 
      -- CP-element group 538: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624__exit__
      -- CP-element group 538: 	 branch_block_stmt_223/ifx_xthen1665_ifx_xend1734
      -- CP-element group 538: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/$exit
      -- CP-element group 538: 	 branch_block_stmt_223/ifx_xthen1665_ifx_xend1734_PhiReq/$entry
      -- CP-element group 538: 	 branch_block_stmt_223/ifx_xthen1665_ifx_xend1734_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_538: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_538"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(532) & zeropad3D_CP_676_elements(537);
      gj_zeropad3D_cp_element_group_538 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(538), clk => clk, reset => reset); --
    end block;
    -- CP-element group 539:  transition  input  bypass 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	523 
    -- CP-element group 539: successors 
    -- CP-element group 539:  members (3) 
      -- CP-element group 539: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_sample_completed_
      -- CP-element group 539: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_Sample/$exit
      -- CP-element group 539: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_Sample/ra
      -- 
    ra_6259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 539_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3630_inst_ack_0, ack => zeropad3D_CP_676_elements(539)); -- 
    -- CP-element group 540:  fork  transition  input  output  bypass 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: 	523 
    -- CP-element group 540: successors 
    -- CP-element group 540: 	541 
    -- CP-element group 540: 	549 
    -- CP-element group 540:  members (9) 
      -- CP-element group 540: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_update_completed_
      -- CP-element group 540: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_Update/$exit
      -- CP-element group 540: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3630_Update/ca
      -- CP-element group 540: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_sample_start_
      -- CP-element group 540: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_Sample/$entry
      -- CP-element group 540: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_Sample/rr
      -- CP-element group 540: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_sample_start_
      -- CP-element group 540: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_Sample/$entry
      -- CP-element group 540: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_Sample/rr
      -- 
    ca_6264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 540_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3630_inst_ack_1, ack => zeropad3D_CP_676_elements(540)); -- 
    rr_6272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(540), ack => type_cast_3694_inst_req_0); -- 
    rr_6382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(540), ack => type_cast_3719_inst_req_0); -- 
    -- CP-element group 541:  transition  input  bypass 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	540 
    -- CP-element group 541: successors 
    -- CP-element group 541:  members (3) 
      -- CP-element group 541: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_sample_completed_
      -- CP-element group 541: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_Sample/$exit
      -- CP-element group 541: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_Sample/ra
      -- 
    ra_6273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 541_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3694_inst_ack_0, ack => zeropad3D_CP_676_elements(541)); -- 
    -- CP-element group 542:  transition  input  output  bypass 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	523 
    -- CP-element group 542: successors 
    -- CP-element group 542: 	543 
    -- CP-element group 542:  members (16) 
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_update_completed_
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_Update/$exit
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3694_Update/ca
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_resized_1
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_scaled_1
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_computed_1
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_resize_1/$entry
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_resize_1/$exit
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_resize_1/index_resize_req
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_resize_1/index_resize_ack
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_scale_1/$entry
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_scale_1/$exit
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_scale_1/scale_rename_req
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_index_scale_1/scale_rename_ack
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_final_index_sum_regn_Sample/$entry
      -- CP-element group 542: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_final_index_sum_regn_Sample/req
      -- 
    ca_6278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 542_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3694_inst_ack_1, ack => zeropad3D_CP_676_elements(542)); -- 
    req_6303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(542), ack => array_obj_ref_3700_index_offset_req_0); -- 
    -- CP-element group 543:  transition  input  bypass 
    -- CP-element group 543: predecessors 
    -- CP-element group 543: 	542 
    -- CP-element group 543: successors 
    -- CP-element group 543: 	558 
    -- CP-element group 543:  members (3) 
      -- CP-element group 543: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_final_index_sum_regn_sample_complete
      -- CP-element group 543: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_final_index_sum_regn_Sample/$exit
      -- CP-element group 543: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_final_index_sum_regn_Sample/ack
      -- 
    ack_6304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 543_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3700_index_offset_ack_0, ack => zeropad3D_CP_676_elements(543)); -- 
    -- CP-element group 544:  transition  input  output  bypass 
    -- CP-element group 544: predecessors 
    -- CP-element group 544: 	523 
    -- CP-element group 544: successors 
    -- CP-element group 544: 	545 
    -- CP-element group 544:  members (11) 
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_sample_start_
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_root_address_calculated
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_offset_calculated
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_final_index_sum_regn_Update/$exit
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_final_index_sum_regn_Update/ack
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_base_plus_offset/$entry
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_base_plus_offset/$exit
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_base_plus_offset/sum_rename_req
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3700_base_plus_offset/sum_rename_ack
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_request/$entry
      -- CP-element group 544: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_request/req
      -- 
    ack_6309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 544_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3700_index_offset_ack_1, ack => zeropad3D_CP_676_elements(544)); -- 
    req_6318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(544), ack => addr_of_3701_final_reg_req_0); -- 
    -- CP-element group 545:  transition  input  bypass 
    -- CP-element group 545: predecessors 
    -- CP-element group 545: 	544 
    -- CP-element group 545: successors 
    -- CP-element group 545:  members (3) 
      -- CP-element group 545: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_sample_completed_
      -- CP-element group 545: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_request/$exit
      -- CP-element group 545: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_request/ack
      -- 
    ack_6319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 545_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3701_final_reg_ack_0, ack => zeropad3D_CP_676_elements(545)); -- 
    -- CP-element group 546:  join  fork  transition  input  output  bypass 
    -- CP-element group 546: predecessors 
    -- CP-element group 546: 	523 
    -- CP-element group 546: successors 
    -- CP-element group 546: 	547 
    -- CP-element group 546:  members (24) 
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_update_completed_
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_complete/$exit
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3701_complete/ack
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_sample_start_
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_base_address_calculated
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_word_address_calculated
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_root_address_calculated
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_base_address_resized
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_base_addr_resize/$entry
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_base_addr_resize/$exit
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_base_addr_resize/base_resize_req
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_base_addr_resize/base_resize_ack
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_base_plus_offset/$entry
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_base_plus_offset/$exit
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_base_plus_offset/sum_rename_req
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_base_plus_offset/sum_rename_ack
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_word_addrgen/$entry
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_word_addrgen/$exit
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_word_addrgen/root_register_req
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_word_addrgen/root_register_ack
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Sample/$entry
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Sample/word_access_start/$entry
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Sample/word_access_start/word_0/$entry
      -- CP-element group 546: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Sample/word_access_start/word_0/rr
      -- 
    ack_6324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 546_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3701_final_reg_ack_1, ack => zeropad3D_CP_676_elements(546)); -- 
    rr_6357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(546), ack => ptr_deref_3705_load_0_req_0); -- 
    -- CP-element group 547:  transition  input  bypass 
    -- CP-element group 547: predecessors 
    -- CP-element group 547: 	546 
    -- CP-element group 547: successors 
    -- CP-element group 547:  members (5) 
      -- CP-element group 547: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_sample_completed_
      -- CP-element group 547: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Sample/$exit
      -- CP-element group 547: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Sample/word_access_start/$exit
      -- CP-element group 547: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Sample/word_access_start/word_0/$exit
      -- CP-element group 547: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Sample/word_access_start/word_0/ra
      -- 
    ra_6358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 547_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3705_load_0_ack_0, ack => zeropad3D_CP_676_elements(547)); -- 
    -- CP-element group 548:  transition  input  bypass 
    -- CP-element group 548: predecessors 
    -- CP-element group 548: 	523 
    -- CP-element group 548: successors 
    -- CP-element group 548: 	555 
    -- CP-element group 548:  members (9) 
      -- CP-element group 548: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_update_completed_
      -- CP-element group 548: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/$exit
      -- CP-element group 548: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/word_access_complete/$exit
      -- CP-element group 548: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/word_access_complete/word_0/$exit
      -- CP-element group 548: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/word_access_complete/word_0/ca
      -- CP-element group 548: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/ptr_deref_3705_Merge/$entry
      -- CP-element group 548: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/ptr_deref_3705_Merge/$exit
      -- CP-element group 548: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/ptr_deref_3705_Merge/merge_req
      -- CP-element group 548: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3705_Update/ptr_deref_3705_Merge/merge_ack
      -- 
    ca_6369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 548_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3705_load_0_ack_1, ack => zeropad3D_CP_676_elements(548)); -- 
    -- CP-element group 549:  transition  input  bypass 
    -- CP-element group 549: predecessors 
    -- CP-element group 549: 	540 
    -- CP-element group 549: successors 
    -- CP-element group 549:  members (3) 
      -- CP-element group 549: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_sample_completed_
      -- CP-element group 549: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_Sample/$exit
      -- CP-element group 549: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_Sample/ra
      -- 
    ra_6383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 549_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3719_inst_ack_0, ack => zeropad3D_CP_676_elements(549)); -- 
    -- CP-element group 550:  transition  input  output  bypass 
    -- CP-element group 550: predecessors 
    -- CP-element group 550: 	523 
    -- CP-element group 550: successors 
    -- CP-element group 550: 	551 
    -- CP-element group 550:  members (16) 
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_update_completed_
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_Update/$exit
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/type_cast_3719_Update/ca
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_resized_1
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_scaled_1
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_computed_1
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_resize_1/$entry
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_resize_1/$exit
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_resize_1/index_resize_req
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_resize_1/index_resize_ack
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_scale_1/$entry
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_scale_1/$exit
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_scale_1/scale_rename_req
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_index_scale_1/scale_rename_ack
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_final_index_sum_regn_Sample/$entry
      -- CP-element group 550: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_final_index_sum_regn_Sample/req
      -- 
    ca_6388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 550_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3719_inst_ack_1, ack => zeropad3D_CP_676_elements(550)); -- 
    req_6413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(550), ack => array_obj_ref_3725_index_offset_req_0); -- 
    -- CP-element group 551:  transition  input  bypass 
    -- CP-element group 551: predecessors 
    -- CP-element group 551: 	550 
    -- CP-element group 551: successors 
    -- CP-element group 551: 	558 
    -- CP-element group 551:  members (3) 
      -- CP-element group 551: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_final_index_sum_regn_sample_complete
      -- CP-element group 551: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_final_index_sum_regn_Sample/$exit
      -- CP-element group 551: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_final_index_sum_regn_Sample/ack
      -- 
    ack_6414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 551_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3725_index_offset_ack_0, ack => zeropad3D_CP_676_elements(551)); -- 
    -- CP-element group 552:  transition  input  output  bypass 
    -- CP-element group 552: predecessors 
    -- CP-element group 552: 	523 
    -- CP-element group 552: successors 
    -- CP-element group 552: 	553 
    -- CP-element group 552:  members (11) 
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_sample_start_
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_root_address_calculated
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_offset_calculated
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_final_index_sum_regn_Update/$exit
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_final_index_sum_regn_Update/ack
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_base_plus_offset/$entry
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_base_plus_offset/$exit
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_base_plus_offset/sum_rename_req
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/array_obj_ref_3725_base_plus_offset/sum_rename_ack
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_request/$entry
      -- CP-element group 552: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_request/req
      -- 
    ack_6419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 552_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3725_index_offset_ack_1, ack => zeropad3D_CP_676_elements(552)); -- 
    req_6428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(552), ack => addr_of_3726_final_reg_req_0); -- 
    -- CP-element group 553:  transition  input  bypass 
    -- CP-element group 553: predecessors 
    -- CP-element group 553: 	552 
    -- CP-element group 553: successors 
    -- CP-element group 553:  members (3) 
      -- CP-element group 553: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_sample_completed_
      -- CP-element group 553: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_request/$exit
      -- CP-element group 553: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_request/ack
      -- 
    ack_6429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 553_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3726_final_reg_ack_0, ack => zeropad3D_CP_676_elements(553)); -- 
    -- CP-element group 554:  fork  transition  input  bypass 
    -- CP-element group 554: predecessors 
    -- CP-element group 554: 	523 
    -- CP-element group 554: successors 
    -- CP-element group 554: 	555 
    -- CP-element group 554:  members (19) 
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_update_completed_
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_complete/$exit
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/addr_of_3726_complete/ack
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_base_address_calculated
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_word_address_calculated
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_root_address_calculated
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_base_address_resized
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_base_addr_resize/$entry
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_base_addr_resize/$exit
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_base_addr_resize/base_resize_req
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_base_addr_resize/base_resize_ack
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_base_plus_offset/$entry
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_base_plus_offset/$exit
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_base_plus_offset/sum_rename_req
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_base_plus_offset/sum_rename_ack
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_word_addrgen/$entry
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_word_addrgen/$exit
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_word_addrgen/root_register_req
      -- CP-element group 554: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_word_addrgen/root_register_ack
      -- 
    ack_6434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 554_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3726_final_reg_ack_1, ack => zeropad3D_CP_676_elements(554)); -- 
    -- CP-element group 555:  join  transition  output  bypass 
    -- CP-element group 555: predecessors 
    -- CP-element group 555: 	548 
    -- CP-element group 555: 	554 
    -- CP-element group 555: successors 
    -- CP-element group 555: 	556 
    -- CP-element group 555:  members (9) 
      -- CP-element group 555: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_sample_start_
      -- CP-element group 555: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/$entry
      -- CP-element group 555: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/ptr_deref_3729_Split/$entry
      -- CP-element group 555: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/ptr_deref_3729_Split/$exit
      -- CP-element group 555: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/ptr_deref_3729_Split/split_req
      -- CP-element group 555: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/ptr_deref_3729_Split/split_ack
      -- CP-element group 555: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/word_access_start/$entry
      -- CP-element group 555: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/word_access_start/word_0/$entry
      -- CP-element group 555: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/word_access_start/word_0/rr
      -- 
    rr_6472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(555), ack => ptr_deref_3729_store_0_req_0); -- 
    zeropad3D_cp_element_group_555: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_555"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(548) & zeropad3D_CP_676_elements(554);
      gj_zeropad3D_cp_element_group_555 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(555), clk => clk, reset => reset); --
    end block;
    -- CP-element group 556:  transition  input  bypass 
    -- CP-element group 556: predecessors 
    -- CP-element group 556: 	555 
    -- CP-element group 556: successors 
    -- CP-element group 556:  members (5) 
      -- CP-element group 556: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_sample_completed_
      -- CP-element group 556: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/$exit
      -- CP-element group 556: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/word_access_start/$exit
      -- CP-element group 556: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/word_access_start/word_0/$exit
      -- CP-element group 556: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Sample/word_access_start/word_0/ra
      -- 
    ra_6473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 556_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3729_store_0_ack_0, ack => zeropad3D_CP_676_elements(556)); -- 
    -- CP-element group 557:  transition  input  bypass 
    -- CP-element group 557: predecessors 
    -- CP-element group 557: 	523 
    -- CP-element group 557: successors 
    -- CP-element group 557: 	558 
    -- CP-element group 557:  members (5) 
      -- CP-element group 557: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_update_completed_
      -- CP-element group 557: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Update/$exit
      -- CP-element group 557: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Update/word_access_complete/$exit
      -- CP-element group 557: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Update/word_access_complete/word_0/$exit
      -- CP-element group 557: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/ptr_deref_3729_Update/word_access_complete/word_0/ca
      -- 
    ca_6484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 557_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3729_store_0_ack_1, ack => zeropad3D_CP_676_elements(557)); -- 
    -- CP-element group 558:  join  transition  place  bypass 
    -- CP-element group 558: predecessors 
    -- CP-element group 558: 	543 
    -- CP-element group 558: 	551 
    -- CP-element group 558: 	557 
    -- CP-element group 558: successors 
    -- CP-element group 558: 	933 
    -- CP-element group 558:  members (5) 
      -- CP-element group 558: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731__exit__
      -- CP-element group 558: 	 branch_block_stmt_223/ifx_xelse1686_ifx_xend1734
      -- CP-element group 558: 	 branch_block_stmt_223/assign_stmt_3631_to_assign_stmt_3731/$exit
      -- CP-element group 558: 	 branch_block_stmt_223/ifx_xelse1686_ifx_xend1734_PhiReq/$entry
      -- CP-element group 558: 	 branch_block_stmt_223/ifx_xelse1686_ifx_xend1734_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_558: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_558"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(543) & zeropad3D_CP_676_elements(551) & zeropad3D_CP_676_elements(557);
      gj_zeropad3D_cp_element_group_558 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(558), clk => clk, reset => reset); --
    end block;
    -- CP-element group 559:  transition  input  bypass 
    -- CP-element group 559: predecessors 
    -- CP-element group 559: 	933 
    -- CP-element group 559: successors 
    -- CP-element group 559:  members (3) 
      -- CP-element group 559: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_sample_completed_
      -- CP-element group 559: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_Sample/$exit
      -- CP-element group 559: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_Sample/ra
      -- 
    ra_6496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 559_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3737_inst_ack_0, ack => zeropad3D_CP_676_elements(559)); -- 
    -- CP-element group 560:  branch  transition  place  input  output  bypass 
    -- CP-element group 560: predecessors 
    -- CP-element group 560: 	933 
    -- CP-element group 560: successors 
    -- CP-element group 560: 	561 
    -- CP-element group 560: 	562 
    -- CP-element group 560:  members (13) 
      -- CP-element group 560: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751__exit__
      -- CP-element group 560: 	 branch_block_stmt_223/if_stmt_3752__entry__
      -- CP-element group 560: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/$exit
      -- CP-element group 560: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_update_completed_
      -- CP-element group 560: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_Update/$exit
      -- CP-element group 560: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_Update/ca
      -- CP-element group 560: 	 branch_block_stmt_223/if_stmt_3752_dead_link/$entry
      -- CP-element group 560: 	 branch_block_stmt_223/if_stmt_3752_eval_test/$entry
      -- CP-element group 560: 	 branch_block_stmt_223/if_stmt_3752_eval_test/$exit
      -- CP-element group 560: 	 branch_block_stmt_223/if_stmt_3752_eval_test/branch_req
      -- CP-element group 560: 	 branch_block_stmt_223/R_cmp1742_3753_place
      -- CP-element group 560: 	 branch_block_stmt_223/if_stmt_3752_if_link/$entry
      -- CP-element group 560: 	 branch_block_stmt_223/if_stmt_3752_else_link/$entry
      -- 
    ca_6501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 560_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3737_inst_ack_1, ack => zeropad3D_CP_676_elements(560)); -- 
    branch_req_6509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(560), ack => if_stmt_3752_branch_req_0); -- 
    -- CP-element group 561:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 561: predecessors 
    -- CP-element group 561: 	560 
    -- CP-element group 561: successors 
    -- CP-element group 561: 	942 
    -- CP-element group 561: 	943 
    -- CP-element group 561: 	945 
    -- CP-element group 561: 	946 
    -- CP-element group 561: 	948 
    -- CP-element group 561: 	949 
    -- CP-element group 561:  members (40) 
      -- CP-element group 561: 	 branch_block_stmt_223/merge_stmt_3758__exit__
      -- CP-element group 561: 	 branch_block_stmt_223/assign_stmt_3764__entry__
      -- CP-element group 561: 	 branch_block_stmt_223/assign_stmt_3764__exit__
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784
      -- CP-element group 561: 	 branch_block_stmt_223/if_stmt_3752_if_link/$exit
      -- CP-element group 561: 	 branch_block_stmt_223/if_stmt_3752_if_link/if_choice_transition
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xend1734_ifx_xthen1744
      -- CP-element group 561: 	 branch_block_stmt_223/assign_stmt_3764/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/assign_stmt_3764/$exit
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xend1734_ifx_xthen1744_PhiReq/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xend1734_ifx_xthen1744_PhiReq/$exit
      -- CP-element group 561: 	 branch_block_stmt_223/merge_stmt_3758_PhiReqMerge
      -- CP-element group 561: 	 branch_block_stmt_223/merge_stmt_3758_PhiAck/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/merge_stmt_3758_PhiAck/$exit
      -- CP-element group 561: 	 branch_block_stmt_223/merge_stmt_3758_PhiAck/dummy
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/SplitProtocol/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/SplitProtocol/Sample/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/SplitProtocol/Sample/rr
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/SplitProtocol/Update/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/SplitProtocol/Update/cr
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/SplitProtocol/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/SplitProtocol/Sample/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/SplitProtocol/Sample/rr
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/SplitProtocol/Update/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/SplitProtocol/Update/cr
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/SplitProtocol/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/SplitProtocol/Sample/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/SplitProtocol/Sample/rr
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/SplitProtocol/Update/$entry
      -- CP-element group 561: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 561_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3752_branch_ack_1, ack => zeropad3D_CP_676_elements(561)); -- 
    rr_9351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(561), ack => type_cast_3821_inst_req_0); -- 
    cr_9356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(561), ack => type_cast_3821_inst_req_1); -- 
    rr_9374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(561), ack => type_cast_3825_inst_req_0); -- 
    cr_9379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(561), ack => type_cast_3825_inst_req_1); -- 
    rr_9397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(561), ack => type_cast_3833_inst_req_0); -- 
    cr_9402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(561), ack => type_cast_3833_inst_req_1); -- 
    -- CP-element group 562:  fork  transition  place  input  output  bypass 
    -- CP-element group 562: predecessors 
    -- CP-element group 562: 	560 
    -- CP-element group 562: successors 
    -- CP-element group 562: 	563 
    -- CP-element group 562: 	564 
    -- CP-element group 562: 	566 
    -- CP-element group 562: 	568 
    -- CP-element group 562:  members (24) 
      -- CP-element group 562: 	 branch_block_stmt_223/merge_stmt_3766__exit__
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807__entry__
      -- CP-element group 562: 	 branch_block_stmt_223/if_stmt_3752_else_link/$exit
      -- CP-element group 562: 	 branch_block_stmt_223/if_stmt_3752_else_link/else_choice_transition
      -- CP-element group 562: 	 branch_block_stmt_223/ifx_xend1734_ifx_xelse1749
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/$entry
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_sample_start_
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_update_start_
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_Sample/$entry
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_Sample/rr
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_Update/$entry
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_Update/cr
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_update_start_
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_Update/$entry
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_Update/cr
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_update_start_
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_Update/$entry
      -- CP-element group 562: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_Update/cr
      -- CP-element group 562: 	 branch_block_stmt_223/ifx_xend1734_ifx_xelse1749_PhiReq/$entry
      -- CP-element group 562: 	 branch_block_stmt_223/ifx_xend1734_ifx_xelse1749_PhiReq/$exit
      -- CP-element group 562: 	 branch_block_stmt_223/merge_stmt_3766_PhiReqMerge
      -- CP-element group 562: 	 branch_block_stmt_223/merge_stmt_3766_PhiAck/$entry
      -- CP-element group 562: 	 branch_block_stmt_223/merge_stmt_3766_PhiAck/$exit
      -- CP-element group 562: 	 branch_block_stmt_223/merge_stmt_3766_PhiAck/dummy
      -- 
    else_choice_transition_6518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 562_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3752_branch_ack_0, ack => zeropad3D_CP_676_elements(562)); -- 
    rr_6534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(562), ack => type_cast_3776_inst_req_0); -- 
    cr_6539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(562), ack => type_cast_3776_inst_req_1); -- 
    cr_6553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(562), ack => type_cast_3785_inst_req_1); -- 
    cr_6567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(562), ack => type_cast_3801_inst_req_1); -- 
    -- CP-element group 563:  transition  input  bypass 
    -- CP-element group 563: predecessors 
    -- CP-element group 563: 	562 
    -- CP-element group 563: successors 
    -- CP-element group 563:  members (3) 
      -- CP-element group 563: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_sample_completed_
      -- CP-element group 563: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_Sample/$exit
      -- CP-element group 563: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_Sample/ra
      -- 
    ra_6535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 563_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3776_inst_ack_0, ack => zeropad3D_CP_676_elements(563)); -- 
    -- CP-element group 564:  transition  input  output  bypass 
    -- CP-element group 564: predecessors 
    -- CP-element group 564: 	562 
    -- CP-element group 564: successors 
    -- CP-element group 564: 	565 
    -- CP-element group 564:  members (6) 
      -- CP-element group 564: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_update_completed_
      -- CP-element group 564: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_Update/$exit
      -- CP-element group 564: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3776_Update/ca
      -- CP-element group 564: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_sample_start_
      -- CP-element group 564: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_Sample/$entry
      -- CP-element group 564: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_Sample/rr
      -- 
    ca_6540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 564_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3776_inst_ack_1, ack => zeropad3D_CP_676_elements(564)); -- 
    rr_6548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(564), ack => type_cast_3785_inst_req_0); -- 
    -- CP-element group 565:  transition  input  bypass 
    -- CP-element group 565: predecessors 
    -- CP-element group 565: 	564 
    -- CP-element group 565: successors 
    -- CP-element group 565:  members (3) 
      -- CP-element group 565: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_sample_completed_
      -- CP-element group 565: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_Sample/$exit
      -- CP-element group 565: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_Sample/ra
      -- 
    ra_6549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 565_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3785_inst_ack_0, ack => zeropad3D_CP_676_elements(565)); -- 
    -- CP-element group 566:  transition  input  output  bypass 
    -- CP-element group 566: predecessors 
    -- CP-element group 566: 	562 
    -- CP-element group 566: successors 
    -- CP-element group 566: 	567 
    -- CP-element group 566:  members (6) 
      -- CP-element group 566: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_update_completed_
      -- CP-element group 566: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_Update/$exit
      -- CP-element group 566: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3785_Update/ca
      -- CP-element group 566: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_sample_start_
      -- CP-element group 566: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_Sample/$entry
      -- CP-element group 566: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_Sample/rr
      -- 
    ca_6554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 566_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3785_inst_ack_1, ack => zeropad3D_CP_676_elements(566)); -- 
    rr_6562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(566), ack => type_cast_3801_inst_req_0); -- 
    -- CP-element group 567:  transition  input  bypass 
    -- CP-element group 567: predecessors 
    -- CP-element group 567: 	566 
    -- CP-element group 567: successors 
    -- CP-element group 567:  members (3) 
      -- CP-element group 567: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_sample_completed_
      -- CP-element group 567: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_Sample/$exit
      -- CP-element group 567: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_Sample/ra
      -- 
    ra_6563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 567_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3801_inst_ack_0, ack => zeropad3D_CP_676_elements(567)); -- 
    -- CP-element group 568:  branch  transition  place  input  output  bypass 
    -- CP-element group 568: predecessors 
    -- CP-element group 568: 	562 
    -- CP-element group 568: successors 
    -- CP-element group 568: 	569 
    -- CP-element group 568: 	570 
    -- CP-element group 568:  members (13) 
      -- CP-element group 568: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807__exit__
      -- CP-element group 568: 	 branch_block_stmt_223/if_stmt_3808__entry__
      -- CP-element group 568: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/$exit
      -- CP-element group 568: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_update_completed_
      -- CP-element group 568: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_Update/$exit
      -- CP-element group 568: 	 branch_block_stmt_223/assign_stmt_3772_to_assign_stmt_3807/type_cast_3801_Update/ca
      -- CP-element group 568: 	 branch_block_stmt_223/if_stmt_3808_dead_link/$entry
      -- CP-element group 568: 	 branch_block_stmt_223/if_stmt_3808_eval_test/$entry
      -- CP-element group 568: 	 branch_block_stmt_223/if_stmt_3808_eval_test/$exit
      -- CP-element group 568: 	 branch_block_stmt_223/if_stmt_3808_eval_test/branch_req
      -- CP-element group 568: 	 branch_block_stmt_223/R_cmp1775_3809_place
      -- CP-element group 568: 	 branch_block_stmt_223/if_stmt_3808_if_link/$entry
      -- CP-element group 568: 	 branch_block_stmt_223/if_stmt_3808_else_link/$entry
      -- 
    ca_6568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 568_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3801_inst_ack_1, ack => zeropad3D_CP_676_elements(568)); -- 
    branch_req_6576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(568), ack => if_stmt_3808_branch_req_0); -- 
    -- CP-element group 569:  fork  transition  place  input  output  bypass 
    -- CP-element group 569: predecessors 
    -- CP-element group 569: 	568 
    -- CP-element group 569: successors 
    -- CP-element group 569: 	571 
    -- CP-element group 569: 	572 
    -- CP-element group 569: 	573 
    -- CP-element group 569: 	574 
    -- CP-element group 569: 	577 
    -- CP-element group 569:  members (27) 
      -- CP-element group 569: 	 branch_block_stmt_223/merge_stmt_3836__exit__
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857__entry__
      -- CP-element group 569: 	 branch_block_stmt_223/if_stmt_3808_if_link/$exit
      -- CP-element group 569: 	 branch_block_stmt_223/if_stmt_3808_if_link/if_choice_transition
      -- CP-element group 569: 	 branch_block_stmt_223/ifx_xelse1749_whilex_xend1785
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/$entry
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_sample_start_
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_update_start_
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_Sample/$entry
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_Sample/rr
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_Update/$entry
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_Update/cr
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_sample_start_
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_update_start_
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_Sample/$entry
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_Sample/rr
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_Update/$entry
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_Update/cr
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_update_start_
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_Update/$entry
      -- CP-element group 569: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_Update/ccr
      -- CP-element group 569: 	 branch_block_stmt_223/ifx_xelse1749_whilex_xend1785_PhiReq/$entry
      -- CP-element group 569: 	 branch_block_stmt_223/ifx_xelse1749_whilex_xend1785_PhiReq/$exit
      -- CP-element group 569: 	 branch_block_stmt_223/merge_stmt_3836_PhiReqMerge
      -- CP-element group 569: 	 branch_block_stmt_223/merge_stmt_3836_PhiAck/$entry
      -- CP-element group 569: 	 branch_block_stmt_223/merge_stmt_3836_PhiAck/$exit
      -- CP-element group 569: 	 branch_block_stmt_223/merge_stmt_3836_PhiAck/dummy
      -- 
    if_choice_transition_6581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 569_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3808_branch_ack_1, ack => zeropad3D_CP_676_elements(569)); -- 
    rr_6598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(569), ack => type_cast_3840_inst_req_0); -- 
    cr_6603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(569), ack => type_cast_3840_inst_req_1); -- 
    rr_6612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(569), ack => type_cast_3844_inst_req_0); -- 
    cr_6617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(569), ack => type_cast_3844_inst_req_1); -- 
    ccr_6631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_6631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(569), ack => call_stmt_3857_call_req_1); -- 
    -- CP-element group 570:  fork  transition  place  input  output  bypass 
    -- CP-element group 570: predecessors 
    -- CP-element group 570: 	568 
    -- CP-element group 570: successors 
    -- CP-element group 570: 	934 
    -- CP-element group 570: 	935 
    -- CP-element group 570: 	936 
    -- CP-element group 570: 	938 
    -- CP-element group 570: 	939 
    -- CP-element group 570:  members (22) 
      -- CP-element group 570: 	 branch_block_stmt_223/if_stmt_3808_else_link/$exit
      -- CP-element group 570: 	 branch_block_stmt_223/if_stmt_3808_else_link/else_choice_transition
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3815/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/SplitProtocol/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/SplitProtocol/Sample/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/SplitProtocol/Sample/rr
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/SplitProtocol/Update/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/SplitProtocol/Update/cr
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/SplitProtocol/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/SplitProtocol/Sample/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/SplitProtocol/Sample/rr
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/SplitProtocol/Update/$entry
      -- CP-element group 570: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 570_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3808_branch_ack_0, ack => zeropad3D_CP_676_elements(570)); -- 
    rr_9302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(570), ack => type_cast_3827_inst_req_0); -- 
    cr_9307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(570), ack => type_cast_3827_inst_req_1); -- 
    rr_9325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(570), ack => type_cast_3831_inst_req_0); -- 
    cr_9330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(570), ack => type_cast_3831_inst_req_1); -- 
    -- CP-element group 571:  transition  input  bypass 
    -- CP-element group 571: predecessors 
    -- CP-element group 571: 	569 
    -- CP-element group 571: successors 
    -- CP-element group 571:  members (3) 
      -- CP-element group 571: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_sample_completed_
      -- CP-element group 571: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_Sample/$exit
      -- CP-element group 571: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_Sample/ra
      -- 
    ra_6599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 571_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3840_inst_ack_0, ack => zeropad3D_CP_676_elements(571)); -- 
    -- CP-element group 572:  transition  input  bypass 
    -- CP-element group 572: predecessors 
    -- CP-element group 572: 	569 
    -- CP-element group 572: successors 
    -- CP-element group 572: 	575 
    -- CP-element group 572:  members (3) 
      -- CP-element group 572: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_update_completed_
      -- CP-element group 572: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_Update/$exit
      -- CP-element group 572: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3840_Update/ca
      -- 
    ca_6604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 572_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3840_inst_ack_1, ack => zeropad3D_CP_676_elements(572)); -- 
    -- CP-element group 573:  transition  input  bypass 
    -- CP-element group 573: predecessors 
    -- CP-element group 573: 	569 
    -- CP-element group 573: successors 
    -- CP-element group 573:  members (3) 
      -- CP-element group 573: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_sample_completed_
      -- CP-element group 573: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_Sample/$exit
      -- CP-element group 573: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_Sample/ra
      -- 
    ra_6613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 573_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3844_inst_ack_0, ack => zeropad3D_CP_676_elements(573)); -- 
    -- CP-element group 574:  transition  input  bypass 
    -- CP-element group 574: predecessors 
    -- CP-element group 574: 	569 
    -- CP-element group 574: successors 
    -- CP-element group 574: 	575 
    -- CP-element group 574:  members (3) 
      -- CP-element group 574: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_update_completed_
      -- CP-element group 574: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_Update/$exit
      -- CP-element group 574: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/type_cast_3844_Update/ca
      -- 
    ca_6618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 574_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3844_inst_ack_1, ack => zeropad3D_CP_676_elements(574)); -- 
    -- CP-element group 575:  join  transition  output  bypass 
    -- CP-element group 575: predecessors 
    -- CP-element group 575: 	572 
    -- CP-element group 575: 	574 
    -- CP-element group 575: successors 
    -- CP-element group 575: 	576 
    -- CP-element group 575:  members (3) 
      -- CP-element group 575: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_sample_start_
      -- CP-element group 575: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_Sample/$entry
      -- CP-element group 575: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_Sample/crr
      -- 
    crr_6626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_6626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(575), ack => call_stmt_3857_call_req_0); -- 
    zeropad3D_cp_element_group_575: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_575"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(572) & zeropad3D_CP_676_elements(574);
      gj_zeropad3D_cp_element_group_575 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(575), clk => clk, reset => reset); --
    end block;
    -- CP-element group 576:  transition  input  bypass 
    -- CP-element group 576: predecessors 
    -- CP-element group 576: 	575 
    -- CP-element group 576: successors 
    -- CP-element group 576:  members (3) 
      -- CP-element group 576: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_sample_completed_
      -- CP-element group 576: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_Sample/$exit
      -- CP-element group 576: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_Sample/cra
      -- 
    cra_6627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 576_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3857_call_ack_0, ack => zeropad3D_CP_676_elements(576)); -- 
    -- CP-element group 577:  transition  place  input  bypass 
    -- CP-element group 577: predecessors 
    -- CP-element group 577: 	569 
    -- CP-element group 577: successors 
    -- CP-element group 577:  members (16) 
      -- CP-element group 577: 	 branch_block_stmt_223/$exit
      -- CP-element group 577: 	 $exit
      -- CP-element group 577: 	 branch_block_stmt_223/branch_block_stmt_223__exit__
      -- CP-element group 577: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857__exit__
      -- CP-element group 577: 	 branch_block_stmt_223/return__
      -- CP-element group 577: 	 branch_block_stmt_223/merge_stmt_3859__exit__
      -- CP-element group 577: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/$exit
      -- CP-element group 577: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_update_completed_
      -- CP-element group 577: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_Update/$exit
      -- CP-element group 577: 	 branch_block_stmt_223/assign_stmt_3841_to_call_stmt_3857/call_stmt_3857_Update/cca
      -- CP-element group 577: 	 branch_block_stmt_223/return___PhiReq/$entry
      -- CP-element group 577: 	 branch_block_stmt_223/return___PhiReq/$exit
      -- CP-element group 577: 	 branch_block_stmt_223/merge_stmt_3859_PhiReqMerge
      -- CP-element group 577: 	 branch_block_stmt_223/merge_stmt_3859_PhiAck/$entry
      -- CP-element group 577: 	 branch_block_stmt_223/merge_stmt_3859_PhiAck/$exit
      -- CP-element group 577: 	 branch_block_stmt_223/merge_stmt_3859_PhiAck/dummy
      -- 
    cca_6632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 577_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3857_call_ack_1, ack => zeropad3D_CP_676_elements(577)); -- 
    -- CP-element group 578:  transition  output  delay-element  bypass 
    -- CP-element group 578: predecessors 
    -- CP-element group 578: 	45 
    -- CP-element group 578: successors 
    -- CP-element group 578: 	582 
    -- CP-element group 578:  members (5) 
      -- CP-element group 578: 	 branch_block_stmt_223/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 578: 	 branch_block_stmt_223/bbx_xnph_forx_xbody_PhiReq/phi_stmt_338/$exit
      -- CP-element group 578: 	 branch_block_stmt_223/bbx_xnph_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/$exit
      -- CP-element group 578: 	 branch_block_stmt_223/bbx_xnph_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_342_konst_delay_trans
      -- CP-element group 578: 	 branch_block_stmt_223/bbx_xnph_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_req
      -- 
    phi_stmt_338_req_6655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_338_req_6655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(578), ack => phi_stmt_338_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(578) is a control-delay.
    cp_element_578_delay: control_delay_element  generic map(name => " 578_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(45), ack => zeropad3D_CP_676_elements(578), clk => clk, reset =>reset);
    -- CP-element group 579:  transition  input  bypass 
    -- CP-element group 579: predecessors 
    -- CP-element group 579: 	87 
    -- CP-element group 579: successors 
    -- CP-element group 579: 	581 
    -- CP-element group 579:  members (2) 
      -- CP-element group 579: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/SplitProtocol/Sample/$exit
      -- CP-element group 579: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/SplitProtocol/Sample/ra
      -- 
    ra_6675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 579_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_344_inst_ack_0, ack => zeropad3D_CP_676_elements(579)); -- 
    -- CP-element group 580:  transition  input  bypass 
    -- CP-element group 580: predecessors 
    -- CP-element group 580: 	87 
    -- CP-element group 580: successors 
    -- CP-element group 580: 	581 
    -- CP-element group 580:  members (2) 
      -- CP-element group 580: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/SplitProtocol/Update/$exit
      -- CP-element group 580: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/SplitProtocol/Update/ca
      -- 
    ca_6680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 580_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_344_inst_ack_1, ack => zeropad3D_CP_676_elements(580)); -- 
    -- CP-element group 581:  join  transition  output  bypass 
    -- CP-element group 581: predecessors 
    -- CP-element group 581: 	579 
    -- CP-element group 581: 	580 
    -- CP-element group 581: successors 
    -- CP-element group 581: 	582 
    -- CP-element group 581:  members (6) 
      -- CP-element group 581: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 581: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/$exit
      -- CP-element group 581: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/$exit
      -- CP-element group 581: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/$exit
      -- CP-element group 581: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_sources/type_cast_344/SplitProtocol/$exit
      -- CP-element group 581: 	 branch_block_stmt_223/forx_xbody_forx_xbody_PhiReq/phi_stmt_338/phi_stmt_338_req
      -- 
    phi_stmt_338_req_6681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_338_req_6681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(581), ack => phi_stmt_338_req_1); -- 
    zeropad3D_cp_element_group_581: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_581"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(579) & zeropad3D_CP_676_elements(580);
      gj_zeropad3D_cp_element_group_581 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(581), clk => clk, reset => reset); --
    end block;
    -- CP-element group 582:  merge  transition  place  bypass 
    -- CP-element group 582: predecessors 
    -- CP-element group 582: 	578 
    -- CP-element group 582: 	581 
    -- CP-element group 582: successors 
    -- CP-element group 582: 	583 
    -- CP-element group 582:  members (2) 
      -- CP-element group 582: 	 branch_block_stmt_223/merge_stmt_337_PhiReqMerge
      -- CP-element group 582: 	 branch_block_stmt_223/merge_stmt_337_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(582) <= OrReduce(zeropad3D_CP_676_elements(578) & zeropad3D_CP_676_elements(581));
    -- CP-element group 583:  fork  transition  place  input  output  bypass 
    -- CP-element group 583: predecessors 
    -- CP-element group 583: 	582 
    -- CP-element group 583: successors 
    -- CP-element group 583: 	73 
    -- CP-element group 583: 	46 
    -- CP-element group 583: 	47 
    -- CP-element group 583: 	49 
    -- CP-element group 583: 	50 
    -- CP-element group 583: 	53 
    -- CP-element group 583: 	57 
    -- CP-element group 583: 	61 
    -- CP-element group 583: 	65 
    -- CP-element group 583: 	69 
    -- CP-element group 583: 	77 
    -- CP-element group 583: 	81 
    -- CP-element group 583: 	84 
    -- CP-element group 583:  members (56) 
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_update_start_
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500__entry__
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_update_start_
      -- CP-element group 583: 	 branch_block_stmt_223/merge_stmt_337__exit__
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_Update/cr
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_update_start_
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_461_Update/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Update/word_access_complete/word_0/cr
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Update/word_access_complete/word_0/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Update/word_access_complete/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_Update/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_Update/cr
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_Update/cr
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/ptr_deref_487_update_start_
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_443_Update/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_update_start_
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_resized_1
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_scaled_1
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_computed_1
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_resize_1/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_resize_1/$exit
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_resize_1/index_resize_req
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_resize_1/index_resize_ack
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_scale_1/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_scale_1/$exit
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_scale_1/scale_rename_req
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_index_scale_1/scale_rename_ack
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_final_index_sum_regn_update_start
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_final_index_sum_regn_Sample/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_final_index_sum_regn_Sample/req
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_final_index_sum_regn_Update/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/array_obj_ref_350_final_index_sum_regn_Update/req
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_complete/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/addr_of_351_complete/req
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_sample_start_
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_Sample/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/RPIPE_zeropad_input_pipe_354_Sample/rr
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_Update/cr
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_update_start_
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_Update/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_358_Update/cr
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_update_start_
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_Update/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_371_Update/cr
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_479_Update/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_update_start_
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_Update/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_389_Update/cr
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_update_start_
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_Update/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_407_Update/cr
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_Update/$entry
      -- CP-element group 583: 	 branch_block_stmt_223/assign_stmt_352_to_assign_stmt_500/type_cast_425_update_start_
      -- CP-element group 583: 	 branch_block_stmt_223/merge_stmt_337_PhiAck/$exit
      -- CP-element group 583: 	 branch_block_stmt_223/merge_stmt_337_PhiAck/phi_stmt_338_ack
      -- 
    phi_stmt_338_ack_6686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 583_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_338_ack_0, ack => zeropad3D_CP_676_elements(583)); -- 
    cr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => type_cast_461_inst_req_1); -- 
    cr_1631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => ptr_deref_487_store_0_req_1); -- 
    cr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => type_cast_425_inst_req_1); -- 
    cr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => type_cast_443_inst_req_1); -- 
    req_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => array_obj_ref_350_index_offset_req_0); -- 
    req_1342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => array_obj_ref_350_index_offset_req_1); -- 
    req_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => addr_of_351_final_reg_req_1); -- 
    rr_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => RPIPE_zeropad_input_pipe_354_inst_req_0); -- 
    cr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => type_cast_479_inst_req_1); -- 
    cr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => type_cast_358_inst_req_1); -- 
    cr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => type_cast_371_inst_req_1); -- 
    cr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => type_cast_389_inst_req_1); -- 
    cr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(583), ack => type_cast_407_inst_req_1); -- 
    -- CP-element group 584:  merge  fork  transition  place  output  bypass 
    -- CP-element group 584: predecessors 
    -- CP-element group 584: 	37 
    -- CP-element group 584: 	86 
    -- CP-element group 584: successors 
    -- CP-element group 584: 	88 
    -- CP-element group 584: 	89 
    -- CP-element group 584: 	90 
    -- CP-element group 584: 	91 
    -- CP-element group 584: 	92 
    -- CP-element group 584: 	93 
    -- CP-element group 584: 	94 
    -- CP-element group 584: 	95 
    -- CP-element group 584: 	96 
    -- CP-element group 584: 	97 
    -- CP-element group 584: 	99 
    -- CP-element group 584: 	100 
    -- CP-element group 584: 	101 
    -- CP-element group 584: 	102 
    -- CP-element group 584: 	103 
    -- CP-element group 584:  members (58) 
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619__entry__
      -- CP-element group 584: 	 branch_block_stmt_223/merge_stmt_509__exit__
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_update_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Sample/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/word_access_complete/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_sample_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Sample/word_access_start/word_0/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_Update/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Sample/word_access_start/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Sample/word_access_start/word_0/rr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_Sample/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_Sample/rr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_sample_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_Update/cr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_Sample/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_update_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_Update/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_root_address_calculated
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_update_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_Update/cr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_word_address_calculated
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_Sample/rr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_update_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_Sample/rr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_Sample/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_update_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_Update/cr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_520_sample_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_Update/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_528_sample_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_Update/cr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_Update/cr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_Sample/rr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_Sample/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_Update/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_update_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_524_Update/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_Sample/rr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_Sample/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_577_sample_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_Update/cr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_Update/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_Sample/rr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_update_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_Sample/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_update_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_516_sample_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_541_sample_start_
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_Update/cr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/type_cast_537_Update/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/word_access_complete/word_0/cr
      -- CP-element group 584: 	 branch_block_stmt_223/assign_stmt_513_to_assign_stmt_619/LOAD_pad_512_Update/word_access_complete/word_0/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/merge_stmt_509_PhiReqMerge
      -- CP-element group 584: 	 branch_block_stmt_223/merge_stmt_509_PhiAck/$entry
      -- CP-element group 584: 	 branch_block_stmt_223/merge_stmt_509_PhiAck/$exit
      -- CP-element group 584: 	 branch_block_stmt_223/merge_stmt_509_PhiAck/dummy
      -- 
    rr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => LOAD_pad_512_load_0_req_0); -- 
    rr_1723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_524_inst_req_0); -- 
    cr_1742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_528_inst_req_1); -- 
    cr_1714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_520_inst_req_1); -- 
    rr_1737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_528_inst_req_0); -- 
    rr_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_520_inst_req_0); -- 
    cr_1784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_577_inst_req_1); -- 
    cr_1700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_516_inst_req_1); -- 
    cr_1728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_524_inst_req_1); -- 
    rr_1779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_577_inst_req_0); -- 
    rr_1695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_516_inst_req_0); -- 
    cr_1770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_541_inst_req_1); -- 
    rr_1765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_541_inst_req_0); -- 
    cr_1756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => type_cast_537_inst_req_1); -- 
    cr_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(584), ack => LOAD_pad_512_load_0_req_1); -- 
    zeropad3D_CP_676_elements(584) <= OrReduce(zeropad3D_CP_676_elements(37) & zeropad3D_CP_676_elements(86));
    -- CP-element group 585:  transition  output  delay-element  bypass 
    -- CP-element group 585: predecessors 
    -- CP-element group 585: 	104 
    -- CP-element group 585: successors 
    -- CP-element group 585: 	588 
    -- CP-element group 585:  members (4) 
      -- CP-element group 585: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_622/$exit
      -- CP-element group 585: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/$exit
      -- CP-element group 585: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_627_konst_delay_trans
      -- CP-element group 585: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_req
      -- 
    phi_stmt_622_req_6720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_622_req_6720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(585), ack => phi_stmt_622_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(585) is a control-delay.
    cp_element_585_delay: control_delay_element  generic map(name => " 585_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(104), ack => zeropad3D_CP_676_elements(585), clk => clk, reset =>reset);
    -- CP-element group 586:  transition  output  delay-element  bypass 
    -- CP-element group 586: predecessors 
    -- CP-element group 586: 	104 
    -- CP-element group 586: successors 
    -- CP-element group 586: 	588 
    -- CP-element group 586:  members (4) 
      -- CP-element group 586: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_630/$exit
      -- CP-element group 586: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/$exit
      -- CP-element group 586: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_634_konst_delay_trans
      -- CP-element group 586: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_req
      -- 
    phi_stmt_630_req_6728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_630_req_6728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(586), ack => phi_stmt_630_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(586) is a control-delay.
    cp_element_586_delay: control_delay_element  generic map(name => " 586_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(104), ack => zeropad3D_CP_676_elements(586), clk => clk, reset =>reset);
    -- CP-element group 587:  transition  output  delay-element  bypass 
    -- CP-element group 587: predecessors 
    -- CP-element group 587: 	104 
    -- CP-element group 587: successors 
    -- CP-element group 587: 	588 
    -- CP-element group 587:  members (4) 
      -- CP-element group 587: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_637/$exit
      -- CP-element group 587: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/$exit
      -- CP-element group 587: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_641_konst_delay_trans
      -- CP-element group 587: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_req
      -- 
    phi_stmt_637_req_6736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_637_req_6736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(587), ack => phi_stmt_637_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(587) is a control-delay.
    cp_element_587_delay: control_delay_element  generic map(name => " 587_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(104), ack => zeropad3D_CP_676_elements(587), clk => clk, reset =>reset);
    -- CP-element group 588:  join  transition  bypass 
    -- CP-element group 588: predecessors 
    -- CP-element group 588: 	585 
    -- CP-element group 588: 	586 
    -- CP-element group 588: 	587 
    -- CP-element group 588: successors 
    -- CP-element group 588: 	599 
    -- CP-element group 588:  members (1) 
      -- CP-element group 588: 	 branch_block_stmt_223/forx_xend_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_588: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_588"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(585) & zeropad3D_CP_676_elements(586) & zeropad3D_CP_676_elements(587);
      gj_zeropad3D_cp_element_group_588 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(588), clk => clk, reset => reset); --
    end block;
    -- CP-element group 589:  transition  input  bypass 
    -- CP-element group 589: predecessors 
    -- CP-element group 589: 	1 
    -- CP-element group 589: successors 
    -- CP-element group 589: 	591 
    -- CP-element group 589:  members (2) 
      -- CP-element group 589: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/SplitProtocol/Sample/$exit
      -- CP-element group 589: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/SplitProtocol/Sample/ra
      -- 
    ra_6756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 589_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_629_inst_ack_0, ack => zeropad3D_CP_676_elements(589)); -- 
    -- CP-element group 590:  transition  input  bypass 
    -- CP-element group 590: predecessors 
    -- CP-element group 590: 	1 
    -- CP-element group 590: successors 
    -- CP-element group 590: 	591 
    -- CP-element group 590:  members (2) 
      -- CP-element group 590: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/SplitProtocol/Update/$exit
      -- CP-element group 590: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/SplitProtocol/Update/ca
      -- 
    ca_6761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 590_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_629_inst_ack_1, ack => zeropad3D_CP_676_elements(590)); -- 
    -- CP-element group 591:  join  transition  output  bypass 
    -- CP-element group 591: predecessors 
    -- CP-element group 591: 	589 
    -- CP-element group 591: 	590 
    -- CP-element group 591: successors 
    -- CP-element group 591: 	598 
    -- CP-element group 591:  members (5) 
      -- CP-element group 591: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/$exit
      -- CP-element group 591: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/$exit
      -- CP-element group 591: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/$exit
      -- CP-element group 591: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_sources/type_cast_629/SplitProtocol/$exit
      -- CP-element group 591: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_622/phi_stmt_622_req
      -- 
    phi_stmt_622_req_6762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_622_req_6762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(591), ack => phi_stmt_622_req_1); -- 
    zeropad3D_cp_element_group_591: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_591"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(589) & zeropad3D_CP_676_elements(590);
      gj_zeropad3D_cp_element_group_591 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(591), clk => clk, reset => reset); --
    end block;
    -- CP-element group 592:  transition  input  bypass 
    -- CP-element group 592: predecessors 
    -- CP-element group 592: 	1 
    -- CP-element group 592: successors 
    -- CP-element group 592: 	594 
    -- CP-element group 592:  members (2) 
      -- CP-element group 592: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/SplitProtocol/Sample/$exit
      -- CP-element group 592: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/SplitProtocol/Sample/ra
      -- 
    ra_6779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 592_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_0, ack => zeropad3D_CP_676_elements(592)); -- 
    -- CP-element group 593:  transition  input  bypass 
    -- CP-element group 593: predecessors 
    -- CP-element group 593: 	1 
    -- CP-element group 593: successors 
    -- CP-element group 593: 	594 
    -- CP-element group 593:  members (2) 
      -- CP-element group 593: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/SplitProtocol/Update/$exit
      -- CP-element group 593: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/SplitProtocol/Update/ca
      -- 
    ca_6784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 593_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_1, ack => zeropad3D_CP_676_elements(593)); -- 
    -- CP-element group 594:  join  transition  output  bypass 
    -- CP-element group 594: predecessors 
    -- CP-element group 594: 	592 
    -- CP-element group 594: 	593 
    -- CP-element group 594: successors 
    -- CP-element group 594: 	598 
    -- CP-element group 594:  members (5) 
      -- CP-element group 594: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/$exit
      -- CP-element group 594: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/$exit
      -- CP-element group 594: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/$exit
      -- CP-element group 594: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_sources/type_cast_636/SplitProtocol/$exit
      -- CP-element group 594: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_630/phi_stmt_630_req
      -- 
    phi_stmt_630_req_6785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_630_req_6785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(594), ack => phi_stmt_630_req_1); -- 
    zeropad3D_cp_element_group_594: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_594"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(592) & zeropad3D_CP_676_elements(593);
      gj_zeropad3D_cp_element_group_594 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(594), clk => clk, reset => reset); --
    end block;
    -- CP-element group 595:  transition  input  bypass 
    -- CP-element group 595: predecessors 
    -- CP-element group 595: 	1 
    -- CP-element group 595: successors 
    -- CP-element group 595: 	597 
    -- CP-element group 595:  members (2) 
      -- CP-element group 595: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/SplitProtocol/Sample/$exit
      -- CP-element group 595: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/SplitProtocol/Sample/ra
      -- 
    ra_6802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 595_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_0, ack => zeropad3D_CP_676_elements(595)); -- 
    -- CP-element group 596:  transition  input  bypass 
    -- CP-element group 596: predecessors 
    -- CP-element group 596: 	1 
    -- CP-element group 596: successors 
    -- CP-element group 596: 	597 
    -- CP-element group 596:  members (2) 
      -- CP-element group 596: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/SplitProtocol/Update/$exit
      -- CP-element group 596: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/SplitProtocol/Update/ca
      -- 
    ca_6807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 596_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_1, ack => zeropad3D_CP_676_elements(596)); -- 
    -- CP-element group 597:  join  transition  output  bypass 
    -- CP-element group 597: predecessors 
    -- CP-element group 597: 	595 
    -- CP-element group 597: 	596 
    -- CP-element group 597: successors 
    -- CP-element group 597: 	598 
    -- CP-element group 597:  members (5) 
      -- CP-element group 597: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/$exit
      -- CP-element group 597: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/$exit
      -- CP-element group 597: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/$exit
      -- CP-element group 597: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_sources/type_cast_643/SplitProtocol/$exit
      -- CP-element group 597: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/phi_stmt_637/phi_stmt_637_req
      -- 
    phi_stmt_637_req_6808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_637_req_6808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(597), ack => phi_stmt_637_req_1); -- 
    zeropad3D_cp_element_group_597: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_597"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(595) & zeropad3D_CP_676_elements(596);
      gj_zeropad3D_cp_element_group_597 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(597), clk => clk, reset => reset); --
    end block;
    -- CP-element group 598:  join  transition  bypass 
    -- CP-element group 598: predecessors 
    -- CP-element group 598: 	591 
    -- CP-element group 598: 	594 
    -- CP-element group 598: 	597 
    -- CP-element group 598: successors 
    -- CP-element group 598: 	599 
    -- CP-element group 598:  members (1) 
      -- CP-element group 598: 	 branch_block_stmt_223/ifx_xend253_whilex_xbody_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_598: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_598"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(591) & zeropad3D_CP_676_elements(594) & zeropad3D_CP_676_elements(597);
      gj_zeropad3D_cp_element_group_598 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(598), clk => clk, reset => reset); --
    end block;
    -- CP-element group 599:  merge  fork  transition  place  bypass 
    -- CP-element group 599: predecessors 
    -- CP-element group 599: 	588 
    -- CP-element group 599: 	598 
    -- CP-element group 599: successors 
    -- CP-element group 599: 	600 
    -- CP-element group 599: 	601 
    -- CP-element group 599: 	602 
    -- CP-element group 599:  members (2) 
      -- CP-element group 599: 	 branch_block_stmt_223/merge_stmt_621_PhiReqMerge
      -- CP-element group 599: 	 branch_block_stmt_223/merge_stmt_621_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(599) <= OrReduce(zeropad3D_CP_676_elements(588) & zeropad3D_CP_676_elements(598));
    -- CP-element group 600:  transition  input  bypass 
    -- CP-element group 600: predecessors 
    -- CP-element group 600: 	599 
    -- CP-element group 600: successors 
    -- CP-element group 600: 	603 
    -- CP-element group 600:  members (1) 
      -- CP-element group 600: 	 branch_block_stmt_223/merge_stmt_621_PhiAck/phi_stmt_622_ack
      -- 
    phi_stmt_622_ack_6813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 600_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_622_ack_0, ack => zeropad3D_CP_676_elements(600)); -- 
    -- CP-element group 601:  transition  input  bypass 
    -- CP-element group 601: predecessors 
    -- CP-element group 601: 	599 
    -- CP-element group 601: successors 
    -- CP-element group 601: 	603 
    -- CP-element group 601:  members (1) 
      -- CP-element group 601: 	 branch_block_stmt_223/merge_stmt_621_PhiAck/phi_stmt_630_ack
      -- 
    phi_stmt_630_ack_6814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 601_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_630_ack_0, ack => zeropad3D_CP_676_elements(601)); -- 
    -- CP-element group 602:  transition  input  bypass 
    -- CP-element group 602: predecessors 
    -- CP-element group 602: 	599 
    -- CP-element group 602: successors 
    -- CP-element group 602: 	603 
    -- CP-element group 602:  members (1) 
      -- CP-element group 602: 	 branch_block_stmt_223/merge_stmt_621_PhiAck/phi_stmt_637_ack
      -- 
    phi_stmt_637_ack_6815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 602_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_637_ack_0, ack => zeropad3D_CP_676_elements(602)); -- 
    -- CP-element group 603:  join  fork  transition  place  output  bypass 
    -- CP-element group 603: predecessors 
    -- CP-element group 603: 	600 
    -- CP-element group 603: 	601 
    -- CP-element group 603: 	602 
    -- CP-element group 603: successors 
    -- CP-element group 603: 	105 
    -- CP-element group 603: 	106 
    -- CP-element group 603:  members (10) 
      -- CP-element group 603: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674__entry__
      -- CP-element group 603: 	 branch_block_stmt_223/merge_stmt_621__exit__
      -- CP-element group 603: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_Update/cr
      -- CP-element group 603: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_Update/$entry
      -- CP-element group 603: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_Sample/rr
      -- CP-element group 603: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_Sample/$entry
      -- CP-element group 603: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_update_start_
      -- CP-element group 603: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/type_cast_648_sample_start_
      -- CP-element group 603: 	 branch_block_stmt_223/assign_stmt_649_to_assign_stmt_674/$entry
      -- CP-element group 603: 	 branch_block_stmt_223/merge_stmt_621_PhiAck/$exit
      -- 
    cr_1801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(603), ack => type_cast_648_inst_req_1); -- 
    rr_1796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(603), ack => type_cast_648_inst_req_0); -- 
    zeropad3D_cp_element_group_603: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_603"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(600) & zeropad3D_CP_676_elements(601) & zeropad3D_CP_676_elements(602);
      gj_zeropad3D_cp_element_group_603 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(603), clk => clk, reset => reset); --
    end block;
    -- CP-element group 604:  merge  fork  transition  place  output  bypass 
    -- CP-element group 604: predecessors 
    -- CP-element group 604: 	108 
    -- CP-element group 604: 	112 
    -- CP-element group 604: successors 
    -- CP-element group 604: 	113 
    -- CP-element group 604: 	114 
    -- CP-element group 604: 	115 
    -- CP-element group 604: 	116 
    -- CP-element group 604: 	119 
    -- CP-element group 604: 	121 
    -- CP-element group 604: 	123 
    -- CP-element group 604: 	125 
    -- CP-element group 604:  members (33) 
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775__entry__
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_update_start_
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_Update/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_sample_start_
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_Sample/rr
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_762_Update/cr
      -- CP-element group 604: 	 branch_block_stmt_223/merge_stmt_718__exit__
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_final_index_sum_regn_update_start
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_update_start_
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_Update/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_complete/req
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_complete/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_Update/cr
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_update_start_
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Update/word_access_complete/word_0/cr
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_Update/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Update/word_access_complete/word_0/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/addr_of_769_update_start_
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_Sample/rr
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_Sample/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_Sample/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Update/word_access_complete/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_update_start_
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/ptr_deref_772_Update/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_727_sample_start_
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_final_index_sum_regn_Update/req
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/array_obj_ref_768_final_index_sum_regn_Update/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/assign_stmt_723_to_assign_stmt_775/type_cast_722_Update/cr
      -- CP-element group 604: 	 branch_block_stmt_223/merge_stmt_718_PhiReqMerge
      -- CP-element group 604: 	 branch_block_stmt_223/merge_stmt_718_PhiAck/$entry
      -- CP-element group 604: 	 branch_block_stmt_223/merge_stmt_718_PhiAck/$exit
      -- CP-element group 604: 	 branch_block_stmt_223/merge_stmt_718_PhiAck/dummy
      -- 
    rr_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(604), ack => type_cast_722_inst_req_0); -- 
    cr_1901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(604), ack => type_cast_762_inst_req_1); -- 
    req_1947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(604), ack => addr_of_769_final_reg_req_1); -- 
    cr_1887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(604), ack => type_cast_727_inst_req_1); -- 
    cr_1997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(604), ack => ptr_deref_772_store_0_req_1); -- 
    rr_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(604), ack => type_cast_727_inst_req_0); -- 
    req_1932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(604), ack => array_obj_ref_768_index_offset_req_1); -- 
    cr_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(604), ack => type_cast_722_inst_req_1); -- 
    zeropad3D_CP_676_elements(604) <= OrReduce(zeropad3D_CP_676_elements(108) & zeropad3D_CP_676_elements(112));
    -- CP-element group 605:  merge  fork  transition  place  output  bypass 
    -- CP-element group 605: predecessors 
    -- CP-element group 605: 	126 
    -- CP-element group 605: 	146 
    -- CP-element group 605: successors 
    -- CP-element group 605: 	147 
    -- CP-element group 605: 	148 
    -- CP-element group 605:  members (13) 
      -- CP-element group 605: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902__entry__
      -- CP-element group 605: 	 branch_block_stmt_223/merge_stmt_884__exit__
      -- CP-element group 605: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/$entry
      -- CP-element group 605: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_sample_start_
      -- CP-element group 605: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_update_start_
      -- CP-element group 605: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_Sample/$entry
      -- CP-element group 605: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_Sample/rr
      -- CP-element group 605: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_Update/$entry
      -- CP-element group 605: 	 branch_block_stmt_223/assign_stmt_889_to_assign_stmt_902/type_cast_888_Update/cr
      -- CP-element group 605: 	 branch_block_stmt_223/merge_stmt_884_PhiReqMerge
      -- CP-element group 605: 	 branch_block_stmt_223/merge_stmt_884_PhiAck/$entry
      -- CP-element group 605: 	 branch_block_stmt_223/merge_stmt_884_PhiAck/$exit
      -- CP-element group 605: 	 branch_block_stmt_223/merge_stmt_884_PhiAck/dummy
      -- 
    rr_2246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(605), ack => type_cast_888_inst_req_0); -- 
    cr_2251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(605), ack => type_cast_888_inst_req_1); -- 
    zeropad3D_CP_676_elements(605) <= OrReduce(zeropad3D_CP_676_elements(126) & zeropad3D_CP_676_elements(146));
    -- CP-element group 606:  transition  input  bypass 
    -- CP-element group 606: predecessors 
    -- CP-element group 606: 	158 
    -- CP-element group 606: successors 
    -- CP-element group 606: 	608 
    -- CP-element group 606:  members (2) 
      -- CP-element group 606: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/SplitProtocol/Sample/$exit
      -- CP-element group 606: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/SplitProtocol/Sample/ra
      -- 
    ra_6905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 606_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_972_inst_ack_0, ack => zeropad3D_CP_676_elements(606)); -- 
    -- CP-element group 607:  transition  input  bypass 
    -- CP-element group 607: predecessors 
    -- CP-element group 607: 	158 
    -- CP-element group 607: successors 
    -- CP-element group 607: 	608 
    -- CP-element group 607:  members (2) 
      -- CP-element group 607: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/SplitProtocol/Update/$exit
      -- CP-element group 607: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/SplitProtocol/Update/ca
      -- 
    ca_6910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 607_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_972_inst_ack_1, ack => zeropad3D_CP_676_elements(607)); -- 
    -- CP-element group 608:  join  transition  output  bypass 
    -- CP-element group 608: predecessors 
    -- CP-element group 608: 	606 
    -- CP-element group 608: 	607 
    -- CP-element group 608: successors 
    -- CP-element group 608: 	613 
    -- CP-element group 608:  members (5) 
      -- CP-element group 608: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/$exit
      -- CP-element group 608: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/$exit
      -- CP-element group 608: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/$exit
      -- CP-element group 608: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_972/SplitProtocol/$exit
      -- CP-element group 608: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_req
      -- 
    phi_stmt_967_req_6911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_967_req_6911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(608), ack => phi_stmt_967_req_1); -- 
    zeropad3D_cp_element_group_608: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_608"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(606) & zeropad3D_CP_676_elements(607);
      gj_zeropad3D_cp_element_group_608 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(608), clk => clk, reset => reset); --
    end block;
    -- CP-element group 609:  transition  input  bypass 
    -- CP-element group 609: predecessors 
    -- CP-element group 609: 	158 
    -- CP-element group 609: successors 
    -- CP-element group 609: 	611 
    -- CP-element group 609:  members (2) 
      -- CP-element group 609: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/SplitProtocol/Sample/ra
      -- CP-element group 609: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/SplitProtocol/Sample/$exit
      -- 
    ra_6928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 609_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_978_inst_ack_0, ack => zeropad3D_CP_676_elements(609)); -- 
    -- CP-element group 610:  transition  input  bypass 
    -- CP-element group 610: predecessors 
    -- CP-element group 610: 	158 
    -- CP-element group 610: successors 
    -- CP-element group 610: 	611 
    -- CP-element group 610:  members (2) 
      -- CP-element group 610: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/SplitProtocol/Update/$exit
      -- CP-element group 610: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/SplitProtocol/Update/ca
      -- 
    ca_6933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 610_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_978_inst_ack_1, ack => zeropad3D_CP_676_elements(610)); -- 
    -- CP-element group 611:  join  transition  output  bypass 
    -- CP-element group 611: predecessors 
    -- CP-element group 611: 	609 
    -- CP-element group 611: 	610 
    -- CP-element group 611: successors 
    -- CP-element group 611: 	613 
    -- CP-element group 611:  members (5) 
      -- CP-element group 611: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_req
      -- CP-element group 611: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/SplitProtocol/$exit
      -- CP-element group 611: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/$exit
      -- CP-element group 611: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/$exit
      -- CP-element group 611: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_978/$exit
      -- 
    phi_stmt_973_req_6934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_973_req_6934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(611), ack => phi_stmt_973_req_1); -- 
    zeropad3D_cp_element_group_611: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_611"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(609) & zeropad3D_CP_676_elements(610);
      gj_zeropad3D_cp_element_group_611 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(611), clk => clk, reset => reset); --
    end block;
    -- CP-element group 612:  transition  output  delay-element  bypass 
    -- CP-element group 612: predecessors 
    -- CP-element group 612: 	158 
    -- CP-element group 612: successors 
    -- CP-element group 612: 	613 
    -- CP-element group 612:  members (4) 
      -- CP-element group 612: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_req
      -- CP-element group 612: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_985_konst_delay_trans
      -- CP-element group 612: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/$exit
      -- CP-element group 612: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/phi_stmt_979/$exit
      -- 
    phi_stmt_979_req_6942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_979_req_6942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(612), ack => phi_stmt_979_req_1); -- 
    -- Element group zeropad3D_CP_676_elements(612) is a control-delay.
    cp_element_612_delay: control_delay_element  generic map(name => " 612_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(158), ack => zeropad3D_CP_676_elements(612), clk => clk, reset =>reset);
    -- CP-element group 613:  join  transition  bypass 
    -- CP-element group 613: predecessors 
    -- CP-element group 613: 	608 
    -- CP-element group 613: 	611 
    -- CP-element group 613: 	612 
    -- CP-element group 613: successors 
    -- CP-element group 613: 	624 
    -- CP-element group 613:  members (1) 
      -- CP-element group 613: 	 branch_block_stmt_223/ifx_xelse217_ifx_xend253_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_613: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_613"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(608) & zeropad3D_CP_676_elements(611) & zeropad3D_CP_676_elements(612);
      gj_zeropad3D_cp_element_group_613 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(613), clk => clk, reset => reset); --
    end block;
    -- CP-element group 614:  transition  input  bypass 
    -- CP-element group 614: predecessors 
    -- CP-element group 614: 	149 
    -- CP-element group 614: successors 
    -- CP-element group 614: 	616 
    -- CP-element group 614:  members (2) 
      -- CP-element group 614: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/SplitProtocol/Sample/$exit
      -- CP-element group 614: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/SplitProtocol/Sample/ra
      -- 
    ra_6962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 614_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_970_inst_ack_0, ack => zeropad3D_CP_676_elements(614)); -- 
    -- CP-element group 615:  transition  input  bypass 
    -- CP-element group 615: predecessors 
    -- CP-element group 615: 	149 
    -- CP-element group 615: successors 
    -- CP-element group 615: 	616 
    -- CP-element group 615:  members (2) 
      -- CP-element group 615: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/SplitProtocol/Update/ca
      -- CP-element group 615: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/SplitProtocol/Update/$exit
      -- 
    ca_6967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 615_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_970_inst_ack_1, ack => zeropad3D_CP_676_elements(615)); -- 
    -- CP-element group 616:  join  transition  output  bypass 
    -- CP-element group 616: predecessors 
    -- CP-element group 616: 	614 
    -- CP-element group 616: 	615 
    -- CP-element group 616: successors 
    -- CP-element group 616: 	623 
    -- CP-element group 616:  members (5) 
      -- CP-element group 616: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/SplitProtocol/$exit
      -- CP-element group 616: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/type_cast_970/$exit
      -- CP-element group 616: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_sources/$exit
      -- CP-element group 616: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/$exit
      -- CP-element group 616: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_967/phi_stmt_967_req
      -- 
    phi_stmt_967_req_6968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_967_req_6968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(616), ack => phi_stmt_967_req_0); -- 
    zeropad3D_cp_element_group_616: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_616"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(614) & zeropad3D_CP_676_elements(615);
      gj_zeropad3D_cp_element_group_616 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(616), clk => clk, reset => reset); --
    end block;
    -- CP-element group 617:  transition  input  bypass 
    -- CP-element group 617: predecessors 
    -- CP-element group 617: 	149 
    -- CP-element group 617: successors 
    -- CP-element group 617: 	619 
    -- CP-element group 617:  members (2) 
      -- CP-element group 617: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/SplitProtocol/Sample/$exit
      -- CP-element group 617: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/SplitProtocol/Sample/ra
      -- 
    ra_6985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 617_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_976_inst_ack_0, ack => zeropad3D_CP_676_elements(617)); -- 
    -- CP-element group 618:  transition  input  bypass 
    -- CP-element group 618: predecessors 
    -- CP-element group 618: 	149 
    -- CP-element group 618: successors 
    -- CP-element group 618: 	619 
    -- CP-element group 618:  members (2) 
      -- CP-element group 618: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/SplitProtocol/Update/$exit
      -- CP-element group 618: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/SplitProtocol/Update/ca
      -- 
    ca_6990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 618_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_976_inst_ack_1, ack => zeropad3D_CP_676_elements(618)); -- 
    -- CP-element group 619:  join  transition  output  bypass 
    -- CP-element group 619: predecessors 
    -- CP-element group 619: 	617 
    -- CP-element group 619: 	618 
    -- CP-element group 619: successors 
    -- CP-element group 619: 	623 
    -- CP-element group 619:  members (5) 
      -- CP-element group 619: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/$exit
      -- CP-element group 619: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/type_cast_976/SplitProtocol/$exit
      -- CP-element group 619: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_sources/$exit
      -- CP-element group 619: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/$exit
      -- CP-element group 619: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_973/phi_stmt_973_req
      -- 
    phi_stmt_973_req_6991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_973_req_6991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(619), ack => phi_stmt_973_req_0); -- 
    zeropad3D_cp_element_group_619: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_619"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(617) & zeropad3D_CP_676_elements(618);
      gj_zeropad3D_cp_element_group_619 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(619), clk => clk, reset => reset); --
    end block;
    -- CP-element group 620:  transition  input  bypass 
    -- CP-element group 620: predecessors 
    -- CP-element group 620: 	149 
    -- CP-element group 620: successors 
    -- CP-element group 620: 	622 
    -- CP-element group 620:  members (2) 
      -- CP-element group 620: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/SplitProtocol/Sample/ra
      -- CP-element group 620: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/SplitProtocol/Sample/$exit
      -- 
    ra_7008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 620_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_982_inst_ack_0, ack => zeropad3D_CP_676_elements(620)); -- 
    -- CP-element group 621:  transition  input  bypass 
    -- CP-element group 621: predecessors 
    -- CP-element group 621: 	149 
    -- CP-element group 621: successors 
    -- CP-element group 621: 	622 
    -- CP-element group 621:  members (2) 
      -- CP-element group 621: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/SplitProtocol/Update/ca
      -- CP-element group 621: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/SplitProtocol/Update/$exit
      -- 
    ca_7013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 621_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_982_inst_ack_1, ack => zeropad3D_CP_676_elements(621)); -- 
    -- CP-element group 622:  join  transition  output  bypass 
    -- CP-element group 622: predecessors 
    -- CP-element group 622: 	620 
    -- CP-element group 622: 	621 
    -- CP-element group 622: successors 
    -- CP-element group 622: 	623 
    -- CP-element group 622:  members (5) 
      -- CP-element group 622: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_req
      -- CP-element group 622: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/SplitProtocol/$exit
      -- CP-element group 622: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/type_cast_982/$exit
      -- CP-element group 622: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/phi_stmt_979_sources/$exit
      -- CP-element group 622: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/phi_stmt_979/$exit
      -- 
    phi_stmt_979_req_7014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_979_req_7014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(622), ack => phi_stmt_979_req_0); -- 
    zeropad3D_cp_element_group_622: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_622"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(620) & zeropad3D_CP_676_elements(621);
      gj_zeropad3D_cp_element_group_622 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(622), clk => clk, reset => reset); --
    end block;
    -- CP-element group 623:  join  transition  bypass 
    -- CP-element group 623: predecessors 
    -- CP-element group 623: 	616 
    -- CP-element group 623: 	619 
    -- CP-element group 623: 	622 
    -- CP-element group 623: successors 
    -- CP-element group 623: 	624 
    -- CP-element group 623:  members (1) 
      -- CP-element group 623: 	 branch_block_stmt_223/ifx_xthen212_ifx_xend253_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_623: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_623"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(616) & zeropad3D_CP_676_elements(619) & zeropad3D_CP_676_elements(622);
      gj_zeropad3D_cp_element_group_623 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(623), clk => clk, reset => reset); --
    end block;
    -- CP-element group 624:  merge  fork  transition  place  bypass 
    -- CP-element group 624: predecessors 
    -- CP-element group 624: 	613 
    -- CP-element group 624: 	623 
    -- CP-element group 624: successors 
    -- CP-element group 624: 	625 
    -- CP-element group 624: 	626 
    -- CP-element group 624: 	627 
    -- CP-element group 624:  members (2) 
      -- CP-element group 624: 	 branch_block_stmt_223/merge_stmt_966_PhiAck/$entry
      -- CP-element group 624: 	 branch_block_stmt_223/merge_stmt_966_PhiReqMerge
      -- 
    zeropad3D_CP_676_elements(624) <= OrReduce(zeropad3D_CP_676_elements(613) & zeropad3D_CP_676_elements(623));
    -- CP-element group 625:  transition  input  bypass 
    -- CP-element group 625: predecessors 
    -- CP-element group 625: 	624 
    -- CP-element group 625: successors 
    -- CP-element group 625: 	628 
    -- CP-element group 625:  members (1) 
      -- CP-element group 625: 	 branch_block_stmt_223/merge_stmt_966_PhiAck/phi_stmt_967_ack
      -- 
    phi_stmt_967_ack_7019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 625_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_967_ack_0, ack => zeropad3D_CP_676_elements(625)); -- 
    -- CP-element group 626:  transition  input  bypass 
    -- CP-element group 626: predecessors 
    -- CP-element group 626: 	624 
    -- CP-element group 626: successors 
    -- CP-element group 626: 	628 
    -- CP-element group 626:  members (1) 
      -- CP-element group 626: 	 branch_block_stmt_223/merge_stmt_966_PhiAck/phi_stmt_973_ack
      -- 
    phi_stmt_973_ack_7020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 626_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_973_ack_0, ack => zeropad3D_CP_676_elements(626)); -- 
    -- CP-element group 627:  transition  input  bypass 
    -- CP-element group 627: predecessors 
    -- CP-element group 627: 	624 
    -- CP-element group 627: successors 
    -- CP-element group 627: 	628 
    -- CP-element group 627:  members (1) 
      -- CP-element group 627: 	 branch_block_stmt_223/merge_stmt_966_PhiAck/phi_stmt_979_ack
      -- 
    phi_stmt_979_ack_7021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 627_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_979_ack_0, ack => zeropad3D_CP_676_elements(627)); -- 
    -- CP-element group 628:  join  transition  bypass 
    -- CP-element group 628: predecessors 
    -- CP-element group 628: 	625 
    -- CP-element group 628: 	626 
    -- CP-element group 628: 	627 
    -- CP-element group 628: successors 
    -- CP-element group 628: 	1 
    -- CP-element group 628:  members (1) 
      -- CP-element group 628: 	 branch_block_stmt_223/merge_stmt_966_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_628: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_628"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(625) & zeropad3D_CP_676_elements(626) & zeropad3D_CP_676_elements(627);
      gj_zeropad3D_cp_element_group_628 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(628), clk => clk, reset => reset); --
    end block;
    -- CP-element group 629:  transition  input  bypass 
    -- CP-element group 629: predecessors 
    -- CP-element group 629: 	2 
    -- CP-element group 629: successors 
    -- CP-element group 629: 	631 
    -- CP-element group 629:  members (2) 
      -- CP-element group 629: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/SplitProtocol/Sample/ra
      -- CP-element group 629: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/SplitProtocol/Sample/$exit
      -- 
    ra_7049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 629_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1039_inst_ack_0, ack => zeropad3D_CP_676_elements(629)); -- 
    -- CP-element group 630:  transition  input  bypass 
    -- CP-element group 630: predecessors 
    -- CP-element group 630: 	2 
    -- CP-element group 630: successors 
    -- CP-element group 630: 	631 
    -- CP-element group 630:  members (2) 
      -- CP-element group 630: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/SplitProtocol/Update/ca
      -- CP-element group 630: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/SplitProtocol/Update/$exit
      -- 
    ca_7054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 630_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1039_inst_ack_1, ack => zeropad3D_CP_676_elements(630)); -- 
    -- CP-element group 631:  join  transition  output  bypass 
    -- CP-element group 631: predecessors 
    -- CP-element group 631: 	629 
    -- CP-element group 631: 	630 
    -- CP-element group 631: successors 
    -- CP-element group 631: 	638 
    -- CP-element group 631:  members (5) 
      -- CP-element group 631: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/$exit
      -- CP-element group 631: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/$exit
      -- CP-element group 631: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_req
      -- CP-element group 631: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/SplitProtocol/$exit
      -- CP-element group 631: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1039/$exit
      -- 
    phi_stmt_1034_req_7055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1034_req_7055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(631), ack => phi_stmt_1034_req_1); -- 
    zeropad3D_cp_element_group_631: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_631"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(629) & zeropad3D_CP_676_elements(630);
      gj_zeropad3D_cp_element_group_631 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(631), clk => clk, reset => reset); --
    end block;
    -- CP-element group 632:  transition  input  bypass 
    -- CP-element group 632: predecessors 
    -- CP-element group 632: 	2 
    -- CP-element group 632: successors 
    -- CP-element group 632: 	634 
    -- CP-element group 632:  members (2) 
      -- CP-element group 632: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/SplitProtocol/Sample/ra
      -- CP-element group 632: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/SplitProtocol/Sample/$exit
      -- 
    ra_7072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 632_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1046_inst_ack_0, ack => zeropad3D_CP_676_elements(632)); -- 
    -- CP-element group 633:  transition  input  bypass 
    -- CP-element group 633: predecessors 
    -- CP-element group 633: 	2 
    -- CP-element group 633: successors 
    -- CP-element group 633: 	634 
    -- CP-element group 633:  members (2) 
      -- CP-element group 633: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/SplitProtocol/Update/ca
      -- CP-element group 633: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/SplitProtocol/Update/$exit
      -- 
    ca_7077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 633_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1046_inst_ack_1, ack => zeropad3D_CP_676_elements(633)); -- 
    -- CP-element group 634:  join  transition  output  bypass 
    -- CP-element group 634: predecessors 
    -- CP-element group 634: 	632 
    -- CP-element group 634: 	633 
    -- CP-element group 634: successors 
    -- CP-element group 634: 	638 
    -- CP-element group 634:  members (5) 
      -- CP-element group 634: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/$exit
      -- CP-element group 634: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/$exit
      -- CP-element group 634: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/$exit
      -- CP-element group 634: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_req
      -- CP-element group 634: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1046/SplitProtocol/$exit
      -- 
    phi_stmt_1040_req_7078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1040_req_7078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(634), ack => phi_stmt_1040_req_1); -- 
    zeropad3D_cp_element_group_634: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_634"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(632) & zeropad3D_CP_676_elements(633);
      gj_zeropad3D_cp_element_group_634 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(634), clk => clk, reset => reset); --
    end block;
    -- CP-element group 635:  transition  input  bypass 
    -- CP-element group 635: predecessors 
    -- CP-element group 635: 	2 
    -- CP-element group 635: successors 
    -- CP-element group 635: 	637 
    -- CP-element group 635:  members (2) 
      -- CP-element group 635: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/SplitProtocol/Sample/ra
      -- CP-element group 635: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/SplitProtocol/Sample/$exit
      -- 
    ra_7095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 635_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1053_inst_ack_0, ack => zeropad3D_CP_676_elements(635)); -- 
    -- CP-element group 636:  transition  input  bypass 
    -- CP-element group 636: predecessors 
    -- CP-element group 636: 	2 
    -- CP-element group 636: successors 
    -- CP-element group 636: 	637 
    -- CP-element group 636:  members (2) 
      -- CP-element group 636: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/SplitProtocol/Update/ca
      -- CP-element group 636: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/SplitProtocol/Update/$exit
      -- 
    ca_7100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 636_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1053_inst_ack_1, ack => zeropad3D_CP_676_elements(636)); -- 
    -- CP-element group 637:  join  transition  output  bypass 
    -- CP-element group 637: predecessors 
    -- CP-element group 637: 	635 
    -- CP-element group 637: 	636 
    -- CP-element group 637: successors 
    -- CP-element group 637: 	638 
    -- CP-element group 637:  members (5) 
      -- CP-element group 637: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_req
      -- CP-element group 637: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/SplitProtocol/$exit
      -- CP-element group 637: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1053/$exit
      -- CP-element group 637: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/$exit
      -- CP-element group 637: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/phi_stmt_1047/$exit
      -- 
    phi_stmt_1047_req_7101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1047_req_7101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(637), ack => phi_stmt_1047_req_1); -- 
    zeropad3D_cp_element_group_637: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_637"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(635) & zeropad3D_CP_676_elements(636);
      gj_zeropad3D_cp_element_group_637 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(637), clk => clk, reset => reset); --
    end block;
    -- CP-element group 638:  join  transition  bypass 
    -- CP-element group 638: predecessors 
    -- CP-element group 638: 	631 
    -- CP-element group 638: 	634 
    -- CP-element group 638: 	637 
    -- CP-element group 638: successors 
    -- CP-element group 638: 	645 
    -- CP-element group 638:  members (1) 
      -- CP-element group 638: 	 branch_block_stmt_223/ifx_xend468_whilex_xbody313_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_638: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_638"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(631) & zeropad3D_CP_676_elements(634) & zeropad3D_CP_676_elements(637);
      gj_zeropad3D_cp_element_group_638 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(638), clk => clk, reset => reset); --
    end block;
    -- CP-element group 639:  transition  input  bypass 
    -- CP-element group 639: predecessors 
    -- CP-element group 639: 	165 
    -- CP-element group 639: successors 
    -- CP-element group 639: 	641 
    -- CP-element group 639:  members (2) 
      -- CP-element group 639: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/SplitProtocol/Sample/$exit
      -- CP-element group 639: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/SplitProtocol/Sample/ra
      -- 
    ra_7121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 639_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1037_inst_ack_0, ack => zeropad3D_CP_676_elements(639)); -- 
    -- CP-element group 640:  transition  input  bypass 
    -- CP-element group 640: predecessors 
    -- CP-element group 640: 	165 
    -- CP-element group 640: successors 
    -- CP-element group 640: 	641 
    -- CP-element group 640:  members (2) 
      -- CP-element group 640: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/SplitProtocol/Update/ca
      -- CP-element group 640: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/SplitProtocol/Update/$exit
      -- 
    ca_7126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 640_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1037_inst_ack_1, ack => zeropad3D_CP_676_elements(640)); -- 
    -- CP-element group 641:  join  transition  output  bypass 
    -- CP-element group 641: predecessors 
    -- CP-element group 641: 	639 
    -- CP-element group 641: 	640 
    -- CP-element group 641: successors 
    -- CP-element group 641: 	644 
    -- CP-element group 641:  members (5) 
      -- CP-element group 641: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/SplitProtocol/$exit
      -- CP-element group 641: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/type_cast_1037/$exit
      -- CP-element group 641: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_sources/$exit
      -- CP-element group 641: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/$exit
      -- CP-element group 641: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1034/phi_stmt_1034_req
      -- 
    phi_stmt_1034_req_7127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1034_req_7127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(641), ack => phi_stmt_1034_req_0); -- 
    zeropad3D_cp_element_group_641: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_641"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(639) & zeropad3D_CP_676_elements(640);
      gj_zeropad3D_cp_element_group_641 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(641), clk => clk, reset => reset); --
    end block;
    -- CP-element group 642:  transition  output  delay-element  bypass 
    -- CP-element group 642: predecessors 
    -- CP-element group 642: 	165 
    -- CP-element group 642: successors 
    -- CP-element group 642: 	644 
    -- CP-element group 642:  members (4) 
      -- CP-element group 642: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_req
      -- CP-element group 642: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/type_cast_1044_konst_delay_trans
      -- CP-element group 642: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1040/phi_stmt_1040_sources/$exit
      -- CP-element group 642: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1040/$exit
      -- 
    phi_stmt_1040_req_7135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1040_req_7135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(642), ack => phi_stmt_1040_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(642) is a control-delay.
    cp_element_642_delay: control_delay_element  generic map(name => " 642_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(165), ack => zeropad3D_CP_676_elements(642), clk => clk, reset =>reset);
    -- CP-element group 643:  transition  output  delay-element  bypass 
    -- CP-element group 643: predecessors 
    -- CP-element group 643: 	165 
    -- CP-element group 643: successors 
    -- CP-element group 643: 	644 
    -- CP-element group 643:  members (4) 
      -- CP-element group 643: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_req
      -- CP-element group 643: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1051_konst_delay_trans
      -- CP-element group 643: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/$exit
      -- CP-element group 643: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/phi_stmt_1047/$exit
      -- 
    phi_stmt_1047_req_7143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1047_req_7143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(643), ack => phi_stmt_1047_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(643) is a control-delay.
    cp_element_643_delay: control_delay_element  generic map(name => " 643_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(165), ack => zeropad3D_CP_676_elements(643), clk => clk, reset =>reset);
    -- CP-element group 644:  join  transition  bypass 
    -- CP-element group 644: predecessors 
    -- CP-element group 644: 	641 
    -- CP-element group 644: 	642 
    -- CP-element group 644: 	643 
    -- CP-element group 644: successors 
    -- CP-element group 644: 	645 
    -- CP-element group 644:  members (1) 
      -- CP-element group 644: 	 branch_block_stmt_223/whilex_xend_whilex_xbody313_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_644: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_644"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(641) & zeropad3D_CP_676_elements(642) & zeropad3D_CP_676_elements(643);
      gj_zeropad3D_cp_element_group_644 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(644), clk => clk, reset => reset); --
    end block;
    -- CP-element group 645:  merge  fork  transition  place  bypass 
    -- CP-element group 645: predecessors 
    -- CP-element group 645: 	638 
    -- CP-element group 645: 	644 
    -- CP-element group 645: successors 
    -- CP-element group 645: 	646 
    -- CP-element group 645: 	647 
    -- CP-element group 645: 	648 
    -- CP-element group 645:  members (2) 
      -- CP-element group 645: 	 branch_block_stmt_223/merge_stmt_1033_PhiAck/$entry
      -- CP-element group 645: 	 branch_block_stmt_223/merge_stmt_1033_PhiReqMerge
      -- 
    zeropad3D_CP_676_elements(645) <= OrReduce(zeropad3D_CP_676_elements(638) & zeropad3D_CP_676_elements(644));
    -- CP-element group 646:  transition  input  bypass 
    -- CP-element group 646: predecessors 
    -- CP-element group 646: 	645 
    -- CP-element group 646: successors 
    -- CP-element group 646: 	649 
    -- CP-element group 646:  members (1) 
      -- CP-element group 646: 	 branch_block_stmt_223/merge_stmt_1033_PhiAck/phi_stmt_1034_ack
      -- 
    phi_stmt_1034_ack_7148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 646_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1034_ack_0, ack => zeropad3D_CP_676_elements(646)); -- 
    -- CP-element group 647:  transition  input  bypass 
    -- CP-element group 647: predecessors 
    -- CP-element group 647: 	645 
    -- CP-element group 647: successors 
    -- CP-element group 647: 	649 
    -- CP-element group 647:  members (1) 
      -- CP-element group 647: 	 branch_block_stmt_223/merge_stmt_1033_PhiAck/phi_stmt_1040_ack
      -- 
    phi_stmt_1040_ack_7149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 647_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1040_ack_0, ack => zeropad3D_CP_676_elements(647)); -- 
    -- CP-element group 648:  transition  input  bypass 
    -- CP-element group 648: predecessors 
    -- CP-element group 648: 	645 
    -- CP-element group 648: successors 
    -- CP-element group 648: 	649 
    -- CP-element group 648:  members (1) 
      -- CP-element group 648: 	 branch_block_stmt_223/merge_stmt_1033_PhiAck/phi_stmt_1047_ack
      -- 
    phi_stmt_1047_ack_7150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 648_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1047_ack_0, ack => zeropad3D_CP_676_elements(648)); -- 
    -- CP-element group 649:  join  fork  transition  place  output  bypass 
    -- CP-element group 649: predecessors 
    -- CP-element group 649: 	646 
    -- CP-element group 649: 	647 
    -- CP-element group 649: 	648 
    -- CP-element group 649: successors 
    -- CP-element group 649: 	166 
    -- CP-element group 649: 	167 
    -- CP-element group 649:  members (10) 
      -- CP-element group 649: 	 branch_block_stmt_223/merge_stmt_1033__exit__
      -- CP-element group 649: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084__entry__
      -- CP-element group 649: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/$entry
      -- CP-element group 649: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_sample_start_
      -- CP-element group 649: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_update_start_
      -- CP-element group 649: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_Sample/$entry
      -- CP-element group 649: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_Sample/rr
      -- CP-element group 649: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_Update/$entry
      -- CP-element group 649: 	 branch_block_stmt_223/assign_stmt_1059_to_assign_stmt_1084/type_cast_1058_Update/cr
      -- CP-element group 649: 	 branch_block_stmt_223/merge_stmt_1033_PhiAck/$exit
      -- 
    rr_2413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(649), ack => type_cast_1058_inst_req_0); -- 
    cr_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(649), ack => type_cast_1058_inst_req_1); -- 
    zeropad3D_cp_element_group_649: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_649"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(646) & zeropad3D_CP_676_elements(647) & zeropad3D_CP_676_elements(648);
      gj_zeropad3D_cp_element_group_649 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(649), clk => clk, reset => reset); --
    end block;
    -- CP-element group 650:  merge  fork  transition  place  output  bypass 
    -- CP-element group 650: predecessors 
    -- CP-element group 650: 	169 
    -- CP-element group 650: 	173 
    -- CP-element group 650: successors 
    -- CP-element group 650: 	174 
    -- CP-element group 650: 	175 
    -- CP-element group 650: 	176 
    -- CP-element group 650: 	177 
    -- CP-element group 650: 	180 
    -- CP-element group 650: 	182 
    -- CP-element group 650: 	184 
    -- CP-element group 650: 	186 
    -- CP-element group 650:  members (33) 
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184__entry__
      -- CP-element group 650: 	 branch_block_stmt_223/merge_stmt_1128__exit__
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_sample_start_
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_update_start_
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_Sample/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_Sample/rr
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_Update/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1132_Update/cr
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_sample_start_
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_update_start_
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_Sample/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_Sample/rr
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_Update/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1137_Update/cr
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_update_start_
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_Update/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/type_cast_1171_Update/cr
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_update_start_
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_final_index_sum_regn_update_start
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_final_index_sum_regn_Update/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/array_obj_ref_1177_final_index_sum_regn_Update/req
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_complete/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/addr_of_1178_complete/req
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_update_start_
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Update/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Update/word_access_complete/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Update/word_access_complete/word_0/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/assign_stmt_1133_to_assign_stmt_1184/ptr_deref_1181_Update/word_access_complete/word_0/cr
      -- CP-element group 650: 	 branch_block_stmt_223/merge_stmt_1128_PhiAck/dummy
      -- CP-element group 650: 	 branch_block_stmt_223/merge_stmt_1128_PhiAck/$exit
      -- CP-element group 650: 	 branch_block_stmt_223/merge_stmt_1128_PhiAck/$entry
      -- CP-element group 650: 	 branch_block_stmt_223/merge_stmt_1128_PhiReqMerge
      -- 
    rr_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(650), ack => type_cast_1132_inst_req_0); -- 
    cr_2490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(650), ack => type_cast_1132_inst_req_1); -- 
    rr_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(650), ack => type_cast_1137_inst_req_0); -- 
    cr_2504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(650), ack => type_cast_1137_inst_req_1); -- 
    cr_2518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(650), ack => type_cast_1171_inst_req_1); -- 
    req_2549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(650), ack => array_obj_ref_1177_index_offset_req_1); -- 
    req_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(650), ack => addr_of_1178_final_reg_req_1); -- 
    cr_2614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(650), ack => ptr_deref_1181_store_0_req_1); -- 
    zeropad3D_CP_676_elements(650) <= OrReduce(zeropad3D_CP_676_elements(169) & zeropad3D_CP_676_elements(173));
    -- CP-element group 651:  merge  fork  transition  place  output  bypass 
    -- CP-element group 651: predecessors 
    -- CP-element group 651: 	187 
    -- CP-element group 651: 	207 
    -- CP-element group 651: successors 
    -- CP-element group 651: 	208 
    -- CP-element group 651: 	209 
    -- CP-element group 651:  members (13) 
      -- CP-element group 651: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311__entry__
      -- CP-element group 651: 	 branch_block_stmt_223/merge_stmt_1293__exit__
      -- CP-element group 651: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_Update/cr
      -- CP-element group 651: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_Update/$entry
      -- CP-element group 651: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_Sample/rr
      -- CP-element group 651: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_Sample/$entry
      -- CP-element group 651: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_update_start_
      -- CP-element group 651: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/type_cast_1297_sample_start_
      -- CP-element group 651: 	 branch_block_stmt_223/assign_stmt_1298_to_assign_stmt_1311/$entry
      -- CP-element group 651: 	 branch_block_stmt_223/merge_stmt_1293_PhiAck/dummy
      -- CP-element group 651: 	 branch_block_stmt_223/merge_stmt_1293_PhiAck/$exit
      -- CP-element group 651: 	 branch_block_stmt_223/merge_stmt_1293_PhiAck/$entry
      -- CP-element group 651: 	 branch_block_stmt_223/merge_stmt_1293_PhiReqMerge
      -- 
    cr_2868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(651), ack => type_cast_1297_inst_req_1); -- 
    rr_2863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(651), ack => type_cast_1297_inst_req_0); -- 
    zeropad3D_CP_676_elements(651) <= OrReduce(zeropad3D_CP_676_elements(187) & zeropad3D_CP_676_elements(207));
    -- CP-element group 652:  transition  input  bypass 
    -- CP-element group 652: predecessors 
    -- CP-element group 652: 	219 
    -- CP-element group 652: successors 
    -- CP-element group 652: 	654 
    -- CP-element group 652:  members (2) 
      -- CP-element group 652: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/SplitProtocol/Sample/ra
      -- CP-element group 652: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/SplitProtocol/Sample/$exit
      -- 
    ra_7240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 652_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_0, ack => zeropad3D_CP_676_elements(652)); -- 
    -- CP-element group 653:  transition  input  bypass 
    -- CP-element group 653: predecessors 
    -- CP-element group 653: 	219 
    -- CP-element group 653: successors 
    -- CP-element group 653: 	654 
    -- CP-element group 653:  members (2) 
      -- CP-element group 653: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/SplitProtocol/Update/$exit
      -- CP-element group 653: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/SplitProtocol/Update/ca
      -- 
    ca_7245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 653_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_1, ack => zeropad3D_CP_676_elements(653)); -- 
    -- CP-element group 654:  join  transition  output  bypass 
    -- CP-element group 654: predecessors 
    -- CP-element group 654: 	652 
    -- CP-element group 654: 	653 
    -- CP-element group 654: successors 
    -- CP-element group 654: 	659 
    -- CP-element group 654:  members (5) 
      -- CP-element group 654: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/SplitProtocol/$exit
      -- CP-element group 654: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1380/$exit
      -- CP-element group 654: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/$exit
      -- CP-element group 654: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_req
      -- CP-element group 654: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1375/$exit
      -- 
    phi_stmt_1375_req_7246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1375_req_7246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(654), ack => phi_stmt_1375_req_1); -- 
    zeropad3D_cp_element_group_654: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_654"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(652) & zeropad3D_CP_676_elements(653);
      gj_zeropad3D_cp_element_group_654 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(654), clk => clk, reset => reset); --
    end block;
    -- CP-element group 655:  transition  input  bypass 
    -- CP-element group 655: predecessors 
    -- CP-element group 655: 	219 
    -- CP-element group 655: successors 
    -- CP-element group 655: 	657 
    -- CP-element group 655:  members (2) 
      -- CP-element group 655: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/SplitProtocol/Sample/ra
      -- CP-element group 655: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/SplitProtocol/Sample/$exit
      -- 
    ra_7263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 655_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_0, ack => zeropad3D_CP_676_elements(655)); -- 
    -- CP-element group 656:  transition  input  bypass 
    -- CP-element group 656: predecessors 
    -- CP-element group 656: 	219 
    -- CP-element group 656: successors 
    -- CP-element group 656: 	657 
    -- CP-element group 656:  members (2) 
      -- CP-element group 656: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/SplitProtocol/Update/ca
      -- CP-element group 656: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/SplitProtocol/Update/$exit
      -- 
    ca_7268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 656_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_1, ack => zeropad3D_CP_676_elements(656)); -- 
    -- CP-element group 657:  join  transition  output  bypass 
    -- CP-element group 657: predecessors 
    -- CP-element group 657: 	655 
    -- CP-element group 657: 	656 
    -- CP-element group 657: successors 
    -- CP-element group 657: 	659 
    -- CP-element group 657:  members (5) 
      -- CP-element group 657: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/$exit
      -- CP-element group 657: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/$exit
      -- CP-element group 657: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/$exit
      -- CP-element group 657: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_req
      -- CP-element group 657: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1386/SplitProtocol/$exit
      -- 
    phi_stmt_1381_req_7269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1381_req_7269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(657), ack => phi_stmt_1381_req_1); -- 
    zeropad3D_cp_element_group_657: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_657"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(655) & zeropad3D_CP_676_elements(656);
      gj_zeropad3D_cp_element_group_657 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(657), clk => clk, reset => reset); --
    end block;
    -- CP-element group 658:  transition  output  delay-element  bypass 
    -- CP-element group 658: predecessors 
    -- CP-element group 658: 	219 
    -- CP-element group 658: successors 
    -- CP-element group 658: 	659 
    -- CP-element group 658:  members (4) 
      -- CP-element group 658: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_req
      -- CP-element group 658: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1393_konst_delay_trans
      -- CP-element group 658: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/$exit
      -- CP-element group 658: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/phi_stmt_1387/$exit
      -- 
    phi_stmt_1387_req_7277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1387_req_7277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(658), ack => phi_stmt_1387_req_1); -- 
    -- Element group zeropad3D_CP_676_elements(658) is a control-delay.
    cp_element_658_delay: control_delay_element  generic map(name => " 658_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(219), ack => zeropad3D_CP_676_elements(658), clk => clk, reset =>reset);
    -- CP-element group 659:  join  transition  bypass 
    -- CP-element group 659: predecessors 
    -- CP-element group 659: 	654 
    -- CP-element group 659: 	657 
    -- CP-element group 659: 	658 
    -- CP-element group 659: successors 
    -- CP-element group 659: 	670 
    -- CP-element group 659:  members (1) 
      -- CP-element group 659: 	 branch_block_stmt_223/ifx_xelse432_ifx_xend468_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_659: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_659"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(654) & zeropad3D_CP_676_elements(657) & zeropad3D_CP_676_elements(658);
      gj_zeropad3D_cp_element_group_659 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(659), clk => clk, reset => reset); --
    end block;
    -- CP-element group 660:  transition  input  bypass 
    -- CP-element group 660: predecessors 
    -- CP-element group 660: 	210 
    -- CP-element group 660: successors 
    -- CP-element group 660: 	662 
    -- CP-element group 660:  members (2) 
      -- CP-element group 660: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/SplitProtocol/Sample/$exit
      -- CP-element group 660: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/SplitProtocol/Sample/ra
      -- 
    ra_7297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 660_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_0, ack => zeropad3D_CP_676_elements(660)); -- 
    -- CP-element group 661:  transition  input  bypass 
    -- CP-element group 661: predecessors 
    -- CP-element group 661: 	210 
    -- CP-element group 661: successors 
    -- CP-element group 661: 	662 
    -- CP-element group 661:  members (2) 
      -- CP-element group 661: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/SplitProtocol/Update/$exit
      -- CP-element group 661: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/SplitProtocol/Update/ca
      -- 
    ca_7302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 661_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_1, ack => zeropad3D_CP_676_elements(661)); -- 
    -- CP-element group 662:  join  transition  output  bypass 
    -- CP-element group 662: predecessors 
    -- CP-element group 662: 	660 
    -- CP-element group 662: 	661 
    -- CP-element group 662: successors 
    -- CP-element group 662: 	669 
    -- CP-element group 662:  members (5) 
      -- CP-element group 662: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/$exit
      -- CP-element group 662: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/$exit
      -- CP-element group 662: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/$exit
      -- CP-element group 662: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_sources/type_cast_1378/SplitProtocol/$exit
      -- CP-element group 662: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1375/phi_stmt_1375_req
      -- 
    phi_stmt_1375_req_7303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1375_req_7303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(662), ack => phi_stmt_1375_req_0); -- 
    zeropad3D_cp_element_group_662: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_662"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(660) & zeropad3D_CP_676_elements(661);
      gj_zeropad3D_cp_element_group_662 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(662), clk => clk, reset => reset); --
    end block;
    -- CP-element group 663:  transition  input  bypass 
    -- CP-element group 663: predecessors 
    -- CP-element group 663: 	210 
    -- CP-element group 663: successors 
    -- CP-element group 663: 	665 
    -- CP-element group 663:  members (2) 
      -- CP-element group 663: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/SplitProtocol/Sample/$exit
      -- CP-element group 663: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/SplitProtocol/Sample/ra
      -- 
    ra_7320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 663_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1384_inst_ack_0, ack => zeropad3D_CP_676_elements(663)); -- 
    -- CP-element group 664:  transition  input  bypass 
    -- CP-element group 664: predecessors 
    -- CP-element group 664: 	210 
    -- CP-element group 664: successors 
    -- CP-element group 664: 	665 
    -- CP-element group 664:  members (2) 
      -- CP-element group 664: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/SplitProtocol/Update/$exit
      -- CP-element group 664: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/SplitProtocol/Update/ca
      -- 
    ca_7325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 664_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1384_inst_ack_1, ack => zeropad3D_CP_676_elements(664)); -- 
    -- CP-element group 665:  join  transition  output  bypass 
    -- CP-element group 665: predecessors 
    -- CP-element group 665: 	663 
    -- CP-element group 665: 	664 
    -- CP-element group 665: successors 
    -- CP-element group 665: 	669 
    -- CP-element group 665:  members (5) 
      -- CP-element group 665: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/$exit
      -- CP-element group 665: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/$exit
      -- CP-element group 665: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/$exit
      -- CP-element group 665: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_sources/type_cast_1384/SplitProtocol/$exit
      -- CP-element group 665: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1381/phi_stmt_1381_req
      -- 
    phi_stmt_1381_req_7326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1381_req_7326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(665), ack => phi_stmt_1381_req_0); -- 
    zeropad3D_cp_element_group_665: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_665"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(663) & zeropad3D_CP_676_elements(664);
      gj_zeropad3D_cp_element_group_665 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(665), clk => clk, reset => reset); --
    end block;
    -- CP-element group 666:  transition  input  bypass 
    -- CP-element group 666: predecessors 
    -- CP-element group 666: 	210 
    -- CP-element group 666: successors 
    -- CP-element group 666: 	668 
    -- CP-element group 666:  members (2) 
      -- CP-element group 666: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/SplitProtocol/Sample/$exit
      -- CP-element group 666: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/SplitProtocol/Sample/ra
      -- 
    ra_7343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 666_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1390_inst_ack_0, ack => zeropad3D_CP_676_elements(666)); -- 
    -- CP-element group 667:  transition  input  bypass 
    -- CP-element group 667: predecessors 
    -- CP-element group 667: 	210 
    -- CP-element group 667: successors 
    -- CP-element group 667: 	668 
    -- CP-element group 667:  members (2) 
      -- CP-element group 667: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/SplitProtocol/Update/$exit
      -- CP-element group 667: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/SplitProtocol/Update/ca
      -- 
    ca_7348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 667_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1390_inst_ack_1, ack => zeropad3D_CP_676_elements(667)); -- 
    -- CP-element group 668:  join  transition  output  bypass 
    -- CP-element group 668: predecessors 
    -- CP-element group 668: 	666 
    -- CP-element group 668: 	667 
    -- CP-element group 668: successors 
    -- CP-element group 668: 	669 
    -- CP-element group 668:  members (5) 
      -- CP-element group 668: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/$exit
      -- CP-element group 668: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/$exit
      -- CP-element group 668: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/$exit
      -- CP-element group 668: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_sources/type_cast_1390/SplitProtocol/$exit
      -- CP-element group 668: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/phi_stmt_1387/phi_stmt_1387_req
      -- 
    phi_stmt_1387_req_7349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1387_req_7349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(668), ack => phi_stmt_1387_req_0); -- 
    zeropad3D_cp_element_group_668: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_668"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(666) & zeropad3D_CP_676_elements(667);
      gj_zeropad3D_cp_element_group_668 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(668), clk => clk, reset => reset); --
    end block;
    -- CP-element group 669:  join  transition  bypass 
    -- CP-element group 669: predecessors 
    -- CP-element group 669: 	662 
    -- CP-element group 669: 	665 
    -- CP-element group 669: 	668 
    -- CP-element group 669: successors 
    -- CP-element group 669: 	670 
    -- CP-element group 669:  members (1) 
      -- CP-element group 669: 	 branch_block_stmt_223/ifx_xthen427_ifx_xend468_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_669: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_669"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(662) & zeropad3D_CP_676_elements(665) & zeropad3D_CP_676_elements(668);
      gj_zeropad3D_cp_element_group_669 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(669), clk => clk, reset => reset); --
    end block;
    -- CP-element group 670:  merge  fork  transition  place  bypass 
    -- CP-element group 670: predecessors 
    -- CP-element group 670: 	659 
    -- CP-element group 670: 	669 
    -- CP-element group 670: successors 
    -- CP-element group 670: 	671 
    -- CP-element group 670: 	672 
    -- CP-element group 670: 	673 
    -- CP-element group 670:  members (2) 
      -- CP-element group 670: 	 branch_block_stmt_223/merge_stmt_1374_PhiReqMerge
      -- CP-element group 670: 	 branch_block_stmt_223/merge_stmt_1374_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(670) <= OrReduce(zeropad3D_CP_676_elements(659) & zeropad3D_CP_676_elements(669));
    -- CP-element group 671:  transition  input  bypass 
    -- CP-element group 671: predecessors 
    -- CP-element group 671: 	670 
    -- CP-element group 671: successors 
    -- CP-element group 671: 	674 
    -- CP-element group 671:  members (1) 
      -- CP-element group 671: 	 branch_block_stmt_223/merge_stmt_1374_PhiAck/phi_stmt_1375_ack
      -- 
    phi_stmt_1375_ack_7354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 671_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1375_ack_0, ack => zeropad3D_CP_676_elements(671)); -- 
    -- CP-element group 672:  transition  input  bypass 
    -- CP-element group 672: predecessors 
    -- CP-element group 672: 	670 
    -- CP-element group 672: successors 
    -- CP-element group 672: 	674 
    -- CP-element group 672:  members (1) 
      -- CP-element group 672: 	 branch_block_stmt_223/merge_stmt_1374_PhiAck/phi_stmt_1381_ack
      -- 
    phi_stmt_1381_ack_7355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 672_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1381_ack_0, ack => zeropad3D_CP_676_elements(672)); -- 
    -- CP-element group 673:  transition  input  bypass 
    -- CP-element group 673: predecessors 
    -- CP-element group 673: 	670 
    -- CP-element group 673: successors 
    -- CP-element group 673: 	674 
    -- CP-element group 673:  members (1) 
      -- CP-element group 673: 	 branch_block_stmt_223/merge_stmt_1374_PhiAck/phi_stmt_1387_ack
      -- 
    phi_stmt_1387_ack_7356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 673_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1387_ack_0, ack => zeropad3D_CP_676_elements(673)); -- 
    -- CP-element group 674:  join  transition  bypass 
    -- CP-element group 674: predecessors 
    -- CP-element group 674: 	671 
    -- CP-element group 674: 	672 
    -- CP-element group 674: 	673 
    -- CP-element group 674: successors 
    -- CP-element group 674: 	2 
    -- CP-element group 674:  members (1) 
      -- CP-element group 674: 	 branch_block_stmt_223/merge_stmt_1374_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_674: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_674"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(671) & zeropad3D_CP_676_elements(672) & zeropad3D_CP_676_elements(673);
      gj_zeropad3D_cp_element_group_674 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(674), clk => clk, reset => reset); --
    end block;
    -- CP-element group 675:  transition  input  bypass 
    -- CP-element group 675: predecessors 
    -- CP-element group 675: 	3 
    -- CP-element group 675: successors 
    -- CP-element group 675: 	677 
    -- CP-element group 675:  members (2) 
      -- CP-element group 675: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/SplitProtocol/Sample/$exit
      -- CP-element group 675: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/SplitProtocol/Sample/ra
      -- 
    ra_7384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 675_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1454_inst_ack_0, ack => zeropad3D_CP_676_elements(675)); -- 
    -- CP-element group 676:  transition  input  bypass 
    -- CP-element group 676: predecessors 
    -- CP-element group 676: 	3 
    -- CP-element group 676: successors 
    -- CP-element group 676: 	677 
    -- CP-element group 676:  members (2) 
      -- CP-element group 676: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/SplitProtocol/Update/$exit
      -- CP-element group 676: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/SplitProtocol/Update/ca
      -- 
    ca_7389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 676_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1454_inst_ack_1, ack => zeropad3D_CP_676_elements(676)); -- 
    -- CP-element group 677:  join  transition  output  bypass 
    -- CP-element group 677: predecessors 
    -- CP-element group 677: 	675 
    -- CP-element group 677: 	676 
    -- CP-element group 677: successors 
    -- CP-element group 677: 	684 
    -- CP-element group 677:  members (5) 
      -- CP-element group 677: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/$exit
      -- CP-element group 677: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/$exit
      -- CP-element group 677: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/$exit
      -- CP-element group 677: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1454/SplitProtocol/$exit
      -- CP-element group 677: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_req
      -- 
    phi_stmt_1448_req_7390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1448_req_7390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(677), ack => phi_stmt_1448_req_1); -- 
    zeropad3D_cp_element_group_677: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_677"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(675) & zeropad3D_CP_676_elements(676);
      gj_zeropad3D_cp_element_group_677 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(677), clk => clk, reset => reset); --
    end block;
    -- CP-element group 678:  transition  input  bypass 
    -- CP-element group 678: predecessors 
    -- CP-element group 678: 	3 
    -- CP-element group 678: successors 
    -- CP-element group 678: 	680 
    -- CP-element group 678:  members (2) 
      -- CP-element group 678: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/SplitProtocol/Sample/$exit
      -- CP-element group 678: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/SplitProtocol/Sample/ra
      -- 
    ra_7407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 678_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1460_inst_ack_0, ack => zeropad3D_CP_676_elements(678)); -- 
    -- CP-element group 679:  transition  input  bypass 
    -- CP-element group 679: predecessors 
    -- CP-element group 679: 	3 
    -- CP-element group 679: successors 
    -- CP-element group 679: 	680 
    -- CP-element group 679:  members (2) 
      -- CP-element group 679: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/SplitProtocol/Update/$exit
      -- CP-element group 679: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/SplitProtocol/Update/ca
      -- 
    ca_7412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 679_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1460_inst_ack_1, ack => zeropad3D_CP_676_elements(679)); -- 
    -- CP-element group 680:  join  transition  output  bypass 
    -- CP-element group 680: predecessors 
    -- CP-element group 680: 	678 
    -- CP-element group 680: 	679 
    -- CP-element group 680: successors 
    -- CP-element group 680: 	684 
    -- CP-element group 680:  members (5) 
      -- CP-element group 680: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/$exit
      -- CP-element group 680: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/$exit
      -- CP-element group 680: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/$exit
      -- CP-element group 680: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1460/SplitProtocol/$exit
      -- CP-element group 680: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_req
      -- 
    phi_stmt_1455_req_7413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1455_req_7413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(680), ack => phi_stmt_1455_req_1); -- 
    zeropad3D_cp_element_group_680: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_680"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(678) & zeropad3D_CP_676_elements(679);
      gj_zeropad3D_cp_element_group_680 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(680), clk => clk, reset => reset); --
    end block;
    -- CP-element group 681:  transition  input  bypass 
    -- CP-element group 681: predecessors 
    -- CP-element group 681: 	3 
    -- CP-element group 681: successors 
    -- CP-element group 681: 	683 
    -- CP-element group 681:  members (2) 
      -- CP-element group 681: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Sample/$exit
      -- CP-element group 681: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Sample/ra
      -- 
    ra_7430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 681_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1467_inst_ack_0, ack => zeropad3D_CP_676_elements(681)); -- 
    -- CP-element group 682:  transition  input  bypass 
    -- CP-element group 682: predecessors 
    -- CP-element group 682: 	3 
    -- CP-element group 682: successors 
    -- CP-element group 682: 	683 
    -- CP-element group 682:  members (2) 
      -- CP-element group 682: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Update/$exit
      -- CP-element group 682: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/Update/ca
      -- 
    ca_7435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 682_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1467_inst_ack_1, ack => zeropad3D_CP_676_elements(682)); -- 
    -- CP-element group 683:  join  transition  output  bypass 
    -- CP-element group 683: predecessors 
    -- CP-element group 683: 	681 
    -- CP-element group 683: 	682 
    -- CP-element group 683: successors 
    -- CP-element group 683: 	684 
    -- CP-element group 683:  members (5) 
      -- CP-element group 683: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/$exit
      -- CP-element group 683: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/$exit
      -- CP-element group 683: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/$exit
      -- CP-element group 683: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1467/SplitProtocol/$exit
      -- CP-element group 683: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_req
      -- 
    phi_stmt_1461_req_7436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1461_req_7436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(683), ack => phi_stmt_1461_req_1); -- 
    zeropad3D_cp_element_group_683: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_683"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(681) & zeropad3D_CP_676_elements(682);
      gj_zeropad3D_cp_element_group_683 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(683), clk => clk, reset => reset); --
    end block;
    -- CP-element group 684:  join  transition  bypass 
    -- CP-element group 684: predecessors 
    -- CP-element group 684: 	677 
    -- CP-element group 684: 	680 
    -- CP-element group 684: 	683 
    -- CP-element group 684: successors 
    -- CP-element group 684: 	691 
    -- CP-element group 684:  members (1) 
      -- CP-element group 684: 	 branch_block_stmt_223/ifx_xend686_whilex_xbody529_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_684: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_684"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(677) & zeropad3D_CP_676_elements(680) & zeropad3D_CP_676_elements(683);
      gj_zeropad3D_cp_element_group_684 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(684), clk => clk, reset => reset); --
    end block;
    -- CP-element group 685:  transition  output  delay-element  bypass 
    -- CP-element group 685: predecessors 
    -- CP-element group 685: 	226 
    -- CP-element group 685: successors 
    -- CP-element group 685: 	690 
    -- CP-element group 685:  members (4) 
      -- CP-element group 685: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1448/$exit
      -- CP-element group 685: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/$exit
      -- CP-element group 685: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_sources/type_cast_1452_konst_delay_trans
      -- CP-element group 685: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1448/phi_stmt_1448_req
      -- 
    phi_stmt_1448_req_7447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1448_req_7447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(685), ack => phi_stmt_1448_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(685) is a control-delay.
    cp_element_685_delay: control_delay_element  generic map(name => " 685_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(226), ack => zeropad3D_CP_676_elements(685), clk => clk, reset =>reset);
    -- CP-element group 686:  transition  input  bypass 
    -- CP-element group 686: predecessors 
    -- CP-element group 686: 	226 
    -- CP-element group 686: successors 
    -- CP-element group 686: 	688 
    -- CP-element group 686:  members (2) 
      -- CP-element group 686: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/SplitProtocol/Sample/$exit
      -- CP-element group 686: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/SplitProtocol/Sample/ra
      -- 
    ra_7464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 686_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1458_inst_ack_0, ack => zeropad3D_CP_676_elements(686)); -- 
    -- CP-element group 687:  transition  input  bypass 
    -- CP-element group 687: predecessors 
    -- CP-element group 687: 	226 
    -- CP-element group 687: successors 
    -- CP-element group 687: 	688 
    -- CP-element group 687:  members (2) 
      -- CP-element group 687: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/SplitProtocol/Update/$exit
      -- CP-element group 687: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/SplitProtocol/Update/ca
      -- 
    ca_7469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 687_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1458_inst_ack_1, ack => zeropad3D_CP_676_elements(687)); -- 
    -- CP-element group 688:  join  transition  output  bypass 
    -- CP-element group 688: predecessors 
    -- CP-element group 688: 	686 
    -- CP-element group 688: 	687 
    -- CP-element group 688: successors 
    -- CP-element group 688: 	690 
    -- CP-element group 688:  members (5) 
      -- CP-element group 688: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/$exit
      -- CP-element group 688: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/$exit
      -- CP-element group 688: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/$exit
      -- CP-element group 688: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_sources/type_cast_1458/SplitProtocol/$exit
      -- CP-element group 688: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1455/phi_stmt_1455_req
      -- 
    phi_stmt_1455_req_7470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1455_req_7470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(688), ack => phi_stmt_1455_req_0); -- 
    zeropad3D_cp_element_group_688: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_688"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(686) & zeropad3D_CP_676_elements(687);
      gj_zeropad3D_cp_element_group_688 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(688), clk => clk, reset => reset); --
    end block;
    -- CP-element group 689:  transition  output  delay-element  bypass 
    -- CP-element group 689: predecessors 
    -- CP-element group 689: 	226 
    -- CP-element group 689: successors 
    -- CP-element group 689: 	690 
    -- CP-element group 689:  members (4) 
      -- CP-element group 689: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1461/$exit
      -- CP-element group 689: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/$exit
      -- CP-element group 689: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_sources/type_cast_1465_konst_delay_trans
      -- CP-element group 689: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/phi_stmt_1461/phi_stmt_1461_req
      -- 
    phi_stmt_1461_req_7478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1461_req_7478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(689), ack => phi_stmt_1461_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(689) is a control-delay.
    cp_element_689_delay: control_delay_element  generic map(name => " 689_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(226), ack => zeropad3D_CP_676_elements(689), clk => clk, reset =>reset);
    -- CP-element group 690:  join  transition  bypass 
    -- CP-element group 690: predecessors 
    -- CP-element group 690: 	685 
    -- CP-element group 690: 	688 
    -- CP-element group 690: 	689 
    -- CP-element group 690: successors 
    -- CP-element group 690: 	691 
    -- CP-element group 690:  members (1) 
      -- CP-element group 690: 	 branch_block_stmt_223/whilex_xend469_whilex_xbody529_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_690: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_690"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(685) & zeropad3D_CP_676_elements(688) & zeropad3D_CP_676_elements(689);
      gj_zeropad3D_cp_element_group_690 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(690), clk => clk, reset => reset); --
    end block;
    -- CP-element group 691:  merge  fork  transition  place  bypass 
    -- CP-element group 691: predecessors 
    -- CP-element group 691: 	684 
    -- CP-element group 691: 	690 
    -- CP-element group 691: successors 
    -- CP-element group 691: 	692 
    -- CP-element group 691: 	693 
    -- CP-element group 691: 	694 
    -- CP-element group 691:  members (2) 
      -- CP-element group 691: 	 branch_block_stmt_223/merge_stmt_1447_PhiReqMerge
      -- CP-element group 691: 	 branch_block_stmt_223/merge_stmt_1447_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(691) <= OrReduce(zeropad3D_CP_676_elements(684) & zeropad3D_CP_676_elements(690));
    -- CP-element group 692:  transition  input  bypass 
    -- CP-element group 692: predecessors 
    -- CP-element group 692: 	691 
    -- CP-element group 692: successors 
    -- CP-element group 692: 	695 
    -- CP-element group 692:  members (1) 
      -- CP-element group 692: 	 branch_block_stmt_223/merge_stmt_1447_PhiAck/phi_stmt_1448_ack
      -- 
    phi_stmt_1448_ack_7483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 692_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1448_ack_0, ack => zeropad3D_CP_676_elements(692)); -- 
    -- CP-element group 693:  transition  input  bypass 
    -- CP-element group 693: predecessors 
    -- CP-element group 693: 	691 
    -- CP-element group 693: successors 
    -- CP-element group 693: 	695 
    -- CP-element group 693:  members (1) 
      -- CP-element group 693: 	 branch_block_stmt_223/merge_stmt_1447_PhiAck/phi_stmt_1455_ack
      -- 
    phi_stmt_1455_ack_7484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 693_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1455_ack_0, ack => zeropad3D_CP_676_elements(693)); -- 
    -- CP-element group 694:  transition  input  bypass 
    -- CP-element group 694: predecessors 
    -- CP-element group 694: 	691 
    -- CP-element group 694: successors 
    -- CP-element group 694: 	695 
    -- CP-element group 694:  members (1) 
      -- CP-element group 694: 	 branch_block_stmt_223/merge_stmt_1447_PhiAck/phi_stmt_1461_ack
      -- 
    phi_stmt_1461_ack_7485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 694_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1461_ack_0, ack => zeropad3D_CP_676_elements(694)); -- 
    -- CP-element group 695:  join  fork  transition  place  output  bypass 
    -- CP-element group 695: predecessors 
    -- CP-element group 695: 	692 
    -- CP-element group 695: 	693 
    -- CP-element group 695: 	694 
    -- CP-element group 695: successors 
    -- CP-element group 695: 	227 
    -- CP-element group 695: 	228 
    -- CP-element group 695:  members (10) 
      -- CP-element group 695: 	 branch_block_stmt_223/merge_stmt_1447__exit__
      -- CP-element group 695: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498__entry__
      -- CP-element group 695: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_Update/cr
      -- CP-element group 695: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_Update/$entry
      -- CP-element group 695: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_Sample/rr
      -- CP-element group 695: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_Sample/$entry
      -- CP-element group 695: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_update_start_
      -- CP-element group 695: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/type_cast_1472_sample_start_
      -- CP-element group 695: 	 branch_block_stmt_223/assign_stmt_1473_to_assign_stmt_1498/$entry
      -- CP-element group 695: 	 branch_block_stmt_223/merge_stmt_1447_PhiAck/$exit
      -- 
    cr_3035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(695), ack => type_cast_1472_inst_req_1); -- 
    rr_3030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(695), ack => type_cast_1472_inst_req_0); -- 
    zeropad3D_cp_element_group_695: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_695"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(692) & zeropad3D_CP_676_elements(693) & zeropad3D_CP_676_elements(694);
      gj_zeropad3D_cp_element_group_695 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(695), clk => clk, reset => reset); --
    end block;
    -- CP-element group 696:  merge  fork  transition  place  output  bypass 
    -- CP-element group 696: predecessors 
    -- CP-element group 696: 	230 
    -- CP-element group 696: 	234 
    -- CP-element group 696: successors 
    -- CP-element group 696: 	235 
    -- CP-element group 696: 	236 
    -- CP-element group 696: 	237 
    -- CP-element group 696: 	238 
    -- CP-element group 696: 	241 
    -- CP-element group 696: 	243 
    -- CP-element group 696: 	245 
    -- CP-element group 696: 	247 
    -- CP-element group 696:  members (33) 
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598__entry__
      -- CP-element group 696: 	 branch_block_stmt_223/merge_stmt_1542__exit__
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_sample_start_
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_update_start_
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_Sample/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_Sample/rr
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_Update/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1546_Update/cr
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_sample_start_
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_update_start_
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_Sample/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_Sample/rr
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_Update/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1551_Update/cr
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_update_start_
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_Update/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/type_cast_1585_Update/cr
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_update_start_
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_final_index_sum_regn_update_start
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_final_index_sum_regn_Update/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/array_obj_ref_1591_final_index_sum_regn_Update/req
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_complete/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/addr_of_1592_complete/req
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_update_start_
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Update/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Update/word_access_complete/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Update/word_access_complete/word_0/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/assign_stmt_1547_to_assign_stmt_1598/ptr_deref_1595_Update/word_access_complete/word_0/cr
      -- CP-element group 696: 	 branch_block_stmt_223/merge_stmt_1542_PhiReqMerge
      -- CP-element group 696: 	 branch_block_stmt_223/merge_stmt_1542_PhiAck/$entry
      -- CP-element group 696: 	 branch_block_stmt_223/merge_stmt_1542_PhiAck/$exit
      -- CP-element group 696: 	 branch_block_stmt_223/merge_stmt_1542_PhiAck/dummy
      -- 
    rr_3102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(696), ack => type_cast_1546_inst_req_0); -- 
    cr_3107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(696), ack => type_cast_1546_inst_req_1); -- 
    rr_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(696), ack => type_cast_1551_inst_req_0); -- 
    cr_3121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(696), ack => type_cast_1551_inst_req_1); -- 
    cr_3135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(696), ack => type_cast_1585_inst_req_1); -- 
    req_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(696), ack => array_obj_ref_1591_index_offset_req_1); -- 
    req_3181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(696), ack => addr_of_1592_final_reg_req_1); -- 
    cr_3231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(696), ack => ptr_deref_1595_store_0_req_1); -- 
    zeropad3D_CP_676_elements(696) <= OrReduce(zeropad3D_CP_676_elements(230) & zeropad3D_CP_676_elements(234));
    -- CP-element group 697:  merge  fork  transition  place  output  bypass 
    -- CP-element group 697: predecessors 
    -- CP-element group 697: 	248 
    -- CP-element group 697: 	268 
    -- CP-element group 697: successors 
    -- CP-element group 697: 	269 
    -- CP-element group 697: 	270 
    -- CP-element group 697:  members (13) 
      -- CP-element group 697: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725__entry__
      -- CP-element group 697: 	 branch_block_stmt_223/merge_stmt_1707__exit__
      -- CP-element group 697: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/$entry
      -- CP-element group 697: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_sample_start_
      -- CP-element group 697: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_update_start_
      -- CP-element group 697: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_Sample/$entry
      -- CP-element group 697: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_Sample/rr
      -- CP-element group 697: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_Update/$entry
      -- CP-element group 697: 	 branch_block_stmt_223/assign_stmt_1712_to_assign_stmt_1725/type_cast_1711_Update/cr
      -- CP-element group 697: 	 branch_block_stmt_223/merge_stmt_1707_PhiReqMerge
      -- CP-element group 697: 	 branch_block_stmt_223/merge_stmt_1707_PhiAck/$entry
      -- CP-element group 697: 	 branch_block_stmt_223/merge_stmt_1707_PhiAck/$exit
      -- CP-element group 697: 	 branch_block_stmt_223/merge_stmt_1707_PhiAck/dummy
      -- 
    rr_3480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(697), ack => type_cast_1711_inst_req_0); -- 
    cr_3485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(697), ack => type_cast_1711_inst_req_1); -- 
    zeropad3D_CP_676_elements(697) <= OrReduce(zeropad3D_CP_676_elements(248) & zeropad3D_CP_676_elements(268));
    -- CP-element group 698:  transition  input  bypass 
    -- CP-element group 698: predecessors 
    -- CP-element group 698: 	280 
    -- CP-element group 698: successors 
    -- CP-element group 698: 	700 
    -- CP-element group 698:  members (2) 
      -- CP-element group 698: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/SplitProtocol/Sample/$exit
      -- CP-element group 698: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/SplitProtocol/Sample/ra
      -- 
    ra_7575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 698_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1808_inst_ack_0, ack => zeropad3D_CP_676_elements(698)); -- 
    -- CP-element group 699:  transition  input  bypass 
    -- CP-element group 699: predecessors 
    -- CP-element group 699: 	280 
    -- CP-element group 699: successors 
    -- CP-element group 699: 	700 
    -- CP-element group 699:  members (2) 
      -- CP-element group 699: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/SplitProtocol/Update/$exit
      -- CP-element group 699: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/SplitProtocol/Update/ca
      -- 
    ca_7580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 699_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1808_inst_ack_1, ack => zeropad3D_CP_676_elements(699)); -- 
    -- CP-element group 700:  join  transition  output  bypass 
    -- CP-element group 700: predecessors 
    -- CP-element group 700: 	698 
    -- CP-element group 700: 	699 
    -- CP-element group 700: successors 
    -- CP-element group 700: 	705 
    -- CP-element group 700:  members (5) 
      -- CP-element group 700: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/$exit
      -- CP-element group 700: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$exit
      -- CP-element group 700: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/$exit
      -- CP-element group 700: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1808/SplitProtocol/$exit
      -- CP-element group 700: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_req
      -- 
    phi_stmt_1803_req_7581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1803_req_7581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(700), ack => phi_stmt_1803_req_1); -- 
    zeropad3D_cp_element_group_700: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_700"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(698) & zeropad3D_CP_676_elements(699);
      gj_zeropad3D_cp_element_group_700 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(700), clk => clk, reset => reset); --
    end block;
    -- CP-element group 701:  transition  input  bypass 
    -- CP-element group 701: predecessors 
    -- CP-element group 701: 	280 
    -- CP-element group 701: successors 
    -- CP-element group 701: 	703 
    -- CP-element group 701:  members (2) 
      -- CP-element group 701: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Sample/$exit
      -- CP-element group 701: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Sample/ra
      -- 
    ra_7598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 701_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1802_inst_ack_0, ack => zeropad3D_CP_676_elements(701)); -- 
    -- CP-element group 702:  transition  input  bypass 
    -- CP-element group 702: predecessors 
    -- CP-element group 702: 	280 
    -- CP-element group 702: successors 
    -- CP-element group 702: 	703 
    -- CP-element group 702:  members (2) 
      -- CP-element group 702: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Update/$exit
      -- CP-element group 702: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/Update/ca
      -- 
    ca_7603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 702_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1802_inst_ack_1, ack => zeropad3D_CP_676_elements(702)); -- 
    -- CP-element group 703:  join  transition  output  bypass 
    -- CP-element group 703: predecessors 
    -- CP-element group 703: 	701 
    -- CP-element group 703: 	702 
    -- CP-element group 703: successors 
    -- CP-element group 703: 	705 
    -- CP-element group 703:  members (5) 
      -- CP-element group 703: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/$exit
      -- CP-element group 703: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/$exit
      -- CP-element group 703: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/$exit
      -- CP-element group 703: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1802/SplitProtocol/$exit
      -- CP-element group 703: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_req
      -- 
    phi_stmt_1797_req_7604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1797_req_7604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(703), ack => phi_stmt_1797_req_1); -- 
    zeropad3D_cp_element_group_703: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_703"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(701) & zeropad3D_CP_676_elements(702);
      gj_zeropad3D_cp_element_group_703 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(703), clk => clk, reset => reset); --
    end block;
    -- CP-element group 704:  transition  output  delay-element  bypass 
    -- CP-element group 704: predecessors 
    -- CP-element group 704: 	280 
    -- CP-element group 704: successors 
    -- CP-element group 704: 	705 
    -- CP-element group 704:  members (4) 
      -- CP-element group 704: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1790/$exit
      -- CP-element group 704: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/$exit
      -- CP-element group 704: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1796_konst_delay_trans
      -- CP-element group 704: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_req
      -- 
    phi_stmt_1790_req_7612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1790_req_7612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(704), ack => phi_stmt_1790_req_1); -- 
    -- Element group zeropad3D_CP_676_elements(704) is a control-delay.
    cp_element_704_delay: control_delay_element  generic map(name => " 704_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(280), ack => zeropad3D_CP_676_elements(704), clk => clk, reset =>reset);
    -- CP-element group 705:  join  transition  bypass 
    -- CP-element group 705: predecessors 
    -- CP-element group 705: 	700 
    -- CP-element group 705: 	703 
    -- CP-element group 705: 	704 
    -- CP-element group 705: successors 
    -- CP-element group 705: 	716 
    -- CP-element group 705:  members (1) 
      -- CP-element group 705: 	 branch_block_stmt_223/ifx_xelse649_ifx_xend686_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_705: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_705"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(700) & zeropad3D_CP_676_elements(703) & zeropad3D_CP_676_elements(704);
      gj_zeropad3D_cp_element_group_705 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(705), clk => clk, reset => reset); --
    end block;
    -- CP-element group 706:  transition  input  bypass 
    -- CP-element group 706: predecessors 
    -- CP-element group 706: 	271 
    -- CP-element group 706: successors 
    -- CP-element group 706: 	708 
    -- CP-element group 706:  members (2) 
      -- CP-element group 706: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/SplitProtocol/Sample/$exit
      -- CP-element group 706: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/SplitProtocol/Sample/ra
      -- 
    ra_7632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 706_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1806_inst_ack_0, ack => zeropad3D_CP_676_elements(706)); -- 
    -- CP-element group 707:  transition  input  bypass 
    -- CP-element group 707: predecessors 
    -- CP-element group 707: 	271 
    -- CP-element group 707: successors 
    -- CP-element group 707: 	708 
    -- CP-element group 707:  members (2) 
      -- CP-element group 707: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/SplitProtocol/Update/$exit
      -- CP-element group 707: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/SplitProtocol/Update/ca
      -- 
    ca_7637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 707_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1806_inst_ack_1, ack => zeropad3D_CP_676_elements(707)); -- 
    -- CP-element group 708:  join  transition  output  bypass 
    -- CP-element group 708: predecessors 
    -- CP-element group 708: 	706 
    -- CP-element group 708: 	707 
    -- CP-element group 708: successors 
    -- CP-element group 708: 	715 
    -- CP-element group 708:  members (5) 
      -- CP-element group 708: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/$exit
      -- CP-element group 708: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$exit
      -- CP-element group 708: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/$exit
      -- CP-element group 708: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1806/SplitProtocol/$exit
      -- CP-element group 708: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1803/phi_stmt_1803_req
      -- 
    phi_stmt_1803_req_7638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1803_req_7638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(708), ack => phi_stmt_1803_req_0); -- 
    zeropad3D_cp_element_group_708: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_708"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(706) & zeropad3D_CP_676_elements(707);
      gj_zeropad3D_cp_element_group_708 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(708), clk => clk, reset => reset); --
    end block;
    -- CP-element group 709:  transition  input  bypass 
    -- CP-element group 709: predecessors 
    -- CP-element group 709: 	271 
    -- CP-element group 709: successors 
    -- CP-element group 709: 	711 
    -- CP-element group 709:  members (2) 
      -- CP-element group 709: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Sample/$exit
      -- CP-element group 709: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Sample/ra
      -- 
    ra_7655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 709_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1800_inst_ack_0, ack => zeropad3D_CP_676_elements(709)); -- 
    -- CP-element group 710:  transition  input  bypass 
    -- CP-element group 710: predecessors 
    -- CP-element group 710: 	271 
    -- CP-element group 710: successors 
    -- CP-element group 710: 	711 
    -- CP-element group 710:  members (2) 
      -- CP-element group 710: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Update/$exit
      -- CP-element group 710: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/Update/ca
      -- 
    ca_7660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 710_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1800_inst_ack_1, ack => zeropad3D_CP_676_elements(710)); -- 
    -- CP-element group 711:  join  transition  output  bypass 
    -- CP-element group 711: predecessors 
    -- CP-element group 711: 	709 
    -- CP-element group 711: 	710 
    -- CP-element group 711: successors 
    -- CP-element group 711: 	715 
    -- CP-element group 711:  members (5) 
      -- CP-element group 711: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/$exit
      -- CP-element group 711: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/$exit
      -- CP-element group 711: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/$exit
      -- CP-element group 711: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_sources/type_cast_1800/SplitProtocol/$exit
      -- CP-element group 711: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1797/phi_stmt_1797_req
      -- 
    phi_stmt_1797_req_7661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1797_req_7661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(711), ack => phi_stmt_1797_req_0); -- 
    zeropad3D_cp_element_group_711: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_711"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(709) & zeropad3D_CP_676_elements(710);
      gj_zeropad3D_cp_element_group_711 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(711), clk => clk, reset => reset); --
    end block;
    -- CP-element group 712:  transition  input  bypass 
    -- CP-element group 712: predecessors 
    -- CP-element group 712: 	271 
    -- CP-element group 712: successors 
    -- CP-element group 712: 	714 
    -- CP-element group 712:  members (2) 
      -- CP-element group 712: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Sample/$exit
      -- CP-element group 712: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Sample/ra
      -- 
    ra_7678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 712_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1793_inst_ack_0, ack => zeropad3D_CP_676_elements(712)); -- 
    -- CP-element group 713:  transition  input  bypass 
    -- CP-element group 713: predecessors 
    -- CP-element group 713: 	271 
    -- CP-element group 713: successors 
    -- CP-element group 713: 	714 
    -- CP-element group 713:  members (2) 
      -- CP-element group 713: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Update/$exit
      -- CP-element group 713: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/Update/ca
      -- 
    ca_7683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 713_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1793_inst_ack_1, ack => zeropad3D_CP_676_elements(713)); -- 
    -- CP-element group 714:  join  transition  output  bypass 
    -- CP-element group 714: predecessors 
    -- CP-element group 714: 	712 
    -- CP-element group 714: 	713 
    -- CP-element group 714: successors 
    -- CP-element group 714: 	715 
    -- CP-element group 714:  members (5) 
      -- CP-element group 714: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/$exit
      -- CP-element group 714: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/$exit
      -- CP-element group 714: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/$exit
      -- CP-element group 714: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_sources/type_cast_1793/SplitProtocol/$exit
      -- CP-element group 714: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/phi_stmt_1790/phi_stmt_1790_req
      -- 
    phi_stmt_1790_req_7684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1790_req_7684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(714), ack => phi_stmt_1790_req_0); -- 
    zeropad3D_cp_element_group_714: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_714"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(712) & zeropad3D_CP_676_elements(713);
      gj_zeropad3D_cp_element_group_714 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(714), clk => clk, reset => reset); --
    end block;
    -- CP-element group 715:  join  transition  bypass 
    -- CP-element group 715: predecessors 
    -- CP-element group 715: 	708 
    -- CP-element group 715: 	711 
    -- CP-element group 715: 	714 
    -- CP-element group 715: successors 
    -- CP-element group 715: 	716 
    -- CP-element group 715:  members (1) 
      -- CP-element group 715: 	 branch_block_stmt_223/ifx_xthen644_ifx_xend686_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_715: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_715"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(708) & zeropad3D_CP_676_elements(711) & zeropad3D_CP_676_elements(714);
      gj_zeropad3D_cp_element_group_715 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(715), clk => clk, reset => reset); --
    end block;
    -- CP-element group 716:  merge  fork  transition  place  bypass 
    -- CP-element group 716: predecessors 
    -- CP-element group 716: 	705 
    -- CP-element group 716: 	715 
    -- CP-element group 716: successors 
    -- CP-element group 716: 	717 
    -- CP-element group 716: 	718 
    -- CP-element group 716: 	719 
    -- CP-element group 716:  members (2) 
      -- CP-element group 716: 	 branch_block_stmt_223/merge_stmt_1789_PhiReqMerge
      -- CP-element group 716: 	 branch_block_stmt_223/merge_stmt_1789_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(716) <= OrReduce(zeropad3D_CP_676_elements(705) & zeropad3D_CP_676_elements(715));
    -- CP-element group 717:  transition  input  bypass 
    -- CP-element group 717: predecessors 
    -- CP-element group 717: 	716 
    -- CP-element group 717: successors 
    -- CP-element group 717: 	720 
    -- CP-element group 717:  members (1) 
      -- CP-element group 717: 	 branch_block_stmt_223/merge_stmt_1789_PhiAck/phi_stmt_1790_ack
      -- 
    phi_stmt_1790_ack_7689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 717_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1790_ack_0, ack => zeropad3D_CP_676_elements(717)); -- 
    -- CP-element group 718:  transition  input  bypass 
    -- CP-element group 718: predecessors 
    -- CP-element group 718: 	716 
    -- CP-element group 718: successors 
    -- CP-element group 718: 	720 
    -- CP-element group 718:  members (1) 
      -- CP-element group 718: 	 branch_block_stmt_223/merge_stmt_1789_PhiAck/phi_stmt_1797_ack
      -- 
    phi_stmt_1797_ack_7690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 718_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1797_ack_0, ack => zeropad3D_CP_676_elements(718)); -- 
    -- CP-element group 719:  transition  input  bypass 
    -- CP-element group 719: predecessors 
    -- CP-element group 719: 	716 
    -- CP-element group 719: successors 
    -- CP-element group 719: 	720 
    -- CP-element group 719:  members (1) 
      -- CP-element group 719: 	 branch_block_stmt_223/merge_stmt_1789_PhiAck/phi_stmt_1803_ack
      -- 
    phi_stmt_1803_ack_7691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 719_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1803_ack_0, ack => zeropad3D_CP_676_elements(719)); -- 
    -- CP-element group 720:  join  transition  bypass 
    -- CP-element group 720: predecessors 
    -- CP-element group 720: 	717 
    -- CP-element group 720: 	718 
    -- CP-element group 720: 	719 
    -- CP-element group 720: successors 
    -- CP-element group 720: 	3 
    -- CP-element group 720:  members (1) 
      -- CP-element group 720: 	 branch_block_stmt_223/merge_stmt_1789_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_720: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_720"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(717) & zeropad3D_CP_676_elements(718) & zeropad3D_CP_676_elements(719);
      gj_zeropad3D_cp_element_group_720 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(720), clk => clk, reset => reset); --
    end block;
    -- CP-element group 721:  transition  input  bypass 
    -- CP-element group 721: predecessors 
    -- CP-element group 721: 	4 
    -- CP-element group 721: successors 
    -- CP-element group 721: 	723 
    -- CP-element group 721:  members (2) 
      -- CP-element group 721: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Sample/$exit
      -- CP-element group 721: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Sample/ra
      -- 
    ra_7719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 721_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1863_inst_ack_0, ack => zeropad3D_CP_676_elements(721)); -- 
    -- CP-element group 722:  transition  input  bypass 
    -- CP-element group 722: predecessors 
    -- CP-element group 722: 	4 
    -- CP-element group 722: successors 
    -- CP-element group 722: 	723 
    -- CP-element group 722:  members (2) 
      -- CP-element group 722: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Update/$exit
      -- CP-element group 722: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Update/ca
      -- 
    ca_7724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 722_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1863_inst_ack_1, ack => zeropad3D_CP_676_elements(722)); -- 
    -- CP-element group 723:  join  transition  output  bypass 
    -- CP-element group 723: predecessors 
    -- CP-element group 723: 	721 
    -- CP-element group 723: 	722 
    -- CP-element group 723: successors 
    -- CP-element group 723: 	730 
    -- CP-element group 723:  members (5) 
      -- CP-element group 723: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/$exit
      -- CP-element group 723: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/$exit
      -- CP-element group 723: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/$exit
      -- CP-element group 723: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/$exit
      -- CP-element group 723: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_req
      -- 
    phi_stmt_1860_req_7725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1860_req_7725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(723), ack => phi_stmt_1860_req_0); -- 
    zeropad3D_cp_element_group_723: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_723"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(721) & zeropad3D_CP_676_elements(722);
      gj_zeropad3D_cp_element_group_723 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(723), clk => clk, reset => reset); --
    end block;
    -- CP-element group 724:  transition  input  bypass 
    -- CP-element group 724: predecessors 
    -- CP-element group 724: 	4 
    -- CP-element group 724: successors 
    -- CP-element group 724: 	726 
    -- CP-element group 724:  members (2) 
      -- CP-element group 724: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Sample/$exit
      -- CP-element group 724: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Sample/ra
      -- 
    ra_7742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 724_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1857_inst_ack_0, ack => zeropad3D_CP_676_elements(724)); -- 
    -- CP-element group 725:  transition  input  bypass 
    -- CP-element group 725: predecessors 
    -- CP-element group 725: 	4 
    -- CP-element group 725: successors 
    -- CP-element group 725: 	726 
    -- CP-element group 725:  members (2) 
      -- CP-element group 725: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Update/$exit
      -- CP-element group 725: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/Update/ca
      -- 
    ca_7747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 725_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1857_inst_ack_1, ack => zeropad3D_CP_676_elements(725)); -- 
    -- CP-element group 726:  join  transition  output  bypass 
    -- CP-element group 726: predecessors 
    -- CP-element group 726: 	724 
    -- CP-element group 726: 	725 
    -- CP-element group 726: successors 
    -- CP-element group 726: 	730 
    -- CP-element group 726:  members (5) 
      -- CP-element group 726: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/$exit
      -- CP-element group 726: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$exit
      -- CP-element group 726: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/$exit
      -- CP-element group 726: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1857/SplitProtocol/$exit
      -- CP-element group 726: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_req
      -- 
    phi_stmt_1854_req_7748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1854_req_7748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(726), ack => phi_stmt_1854_req_0); -- 
    zeropad3D_cp_element_group_726: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_726"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(724) & zeropad3D_CP_676_elements(725);
      gj_zeropad3D_cp_element_group_726 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(726), clk => clk, reset => reset); --
    end block;
    -- CP-element group 727:  transition  input  bypass 
    -- CP-element group 727: predecessors 
    -- CP-element group 727: 	4 
    -- CP-element group 727: successors 
    -- CP-element group 727: 	729 
    -- CP-element group 727:  members (2) 
      -- CP-element group 727: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/SplitProtocol/Sample/$exit
      -- CP-element group 727: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/SplitProtocol/Sample/ra
      -- 
    ra_7765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 727_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1850_inst_ack_0, ack => zeropad3D_CP_676_elements(727)); -- 
    -- CP-element group 728:  transition  input  bypass 
    -- CP-element group 728: predecessors 
    -- CP-element group 728: 	4 
    -- CP-element group 728: successors 
    -- CP-element group 728: 	729 
    -- CP-element group 728:  members (2) 
      -- CP-element group 728: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/SplitProtocol/Update/$exit
      -- CP-element group 728: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/SplitProtocol/Update/ca
      -- 
    ca_7770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 728_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1850_inst_ack_1, ack => zeropad3D_CP_676_elements(728)); -- 
    -- CP-element group 729:  join  transition  output  bypass 
    -- CP-element group 729: predecessors 
    -- CP-element group 729: 	727 
    -- CP-element group 729: 	728 
    -- CP-element group 729: successors 
    -- CP-element group 729: 	730 
    -- CP-element group 729:  members (5) 
      -- CP-element group 729: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/$exit
      -- CP-element group 729: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/$exit
      -- CP-element group 729: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/$exit
      -- CP-element group 729: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1850/SplitProtocol/$exit
      -- CP-element group 729: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_req
      -- 
    phi_stmt_1847_req_7771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1847_req_7771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(729), ack => phi_stmt_1847_req_0); -- 
    zeropad3D_cp_element_group_729: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_729"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(727) & zeropad3D_CP_676_elements(728);
      gj_zeropad3D_cp_element_group_729 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(729), clk => clk, reset => reset); --
    end block;
    -- CP-element group 730:  join  transition  bypass 
    -- CP-element group 730: predecessors 
    -- CP-element group 730: 	723 
    -- CP-element group 730: 	726 
    -- CP-element group 730: 	729 
    -- CP-element group 730: successors 
    -- CP-element group 730: 	739 
    -- CP-element group 730:  members (1) 
      -- CP-element group 730: 	 branch_block_stmt_223/ifx_xend906_whilex_xbody751_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_730: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_730"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(723) & zeropad3D_CP_676_elements(726) & zeropad3D_CP_676_elements(729);
      gj_zeropad3D_cp_element_group_730 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(730), clk => clk, reset => reset); --
    end block;
    -- CP-element group 731:  transition  input  bypass 
    -- CP-element group 731: predecessors 
    -- CP-element group 731: 	284 
    -- CP-element group 731: successors 
    -- CP-element group 731: 	733 
    -- CP-element group 731:  members (2) 
      -- CP-element group 731: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/SplitProtocol/Sample/$exit
      -- CP-element group 731: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/SplitProtocol/Sample/ra
      -- 
    ra_7791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 731_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1865_inst_ack_0, ack => zeropad3D_CP_676_elements(731)); -- 
    -- CP-element group 732:  transition  input  bypass 
    -- CP-element group 732: predecessors 
    -- CP-element group 732: 	284 
    -- CP-element group 732: successors 
    -- CP-element group 732: 	733 
    -- CP-element group 732:  members (2) 
      -- CP-element group 732: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/SplitProtocol/Update/$exit
      -- CP-element group 732: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/SplitProtocol/Update/ca
      -- 
    ca_7796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 732_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1865_inst_ack_1, ack => zeropad3D_CP_676_elements(732)); -- 
    -- CP-element group 733:  join  transition  output  bypass 
    -- CP-element group 733: predecessors 
    -- CP-element group 733: 	731 
    -- CP-element group 733: 	732 
    -- CP-element group 733: successors 
    -- CP-element group 733: 	738 
    -- CP-element group 733:  members (5) 
      -- CP-element group 733: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/$exit
      -- CP-element group 733: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/$exit
      -- CP-element group 733: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/$exit
      -- CP-element group 733: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1865/SplitProtocol/$exit
      -- CP-element group 733: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1860/phi_stmt_1860_req
      -- 
    phi_stmt_1860_req_7797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1860_req_7797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(733), ack => phi_stmt_1860_req_1); -- 
    zeropad3D_cp_element_group_733: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_733"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(731) & zeropad3D_CP_676_elements(732);
      gj_zeropad3D_cp_element_group_733 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(733), clk => clk, reset => reset); --
    end block;
    -- CP-element group 734:  transition  input  bypass 
    -- CP-element group 734: predecessors 
    -- CP-element group 734: 	284 
    -- CP-element group 734: successors 
    -- CP-element group 734: 	736 
    -- CP-element group 734:  members (2) 
      -- CP-element group 734: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/SplitProtocol/Sample/$exit
      -- CP-element group 734: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/SplitProtocol/Sample/ra
      -- 
    ra_7814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 734_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1859_inst_ack_0, ack => zeropad3D_CP_676_elements(734)); -- 
    -- CP-element group 735:  transition  input  bypass 
    -- CP-element group 735: predecessors 
    -- CP-element group 735: 	284 
    -- CP-element group 735: successors 
    -- CP-element group 735: 	736 
    -- CP-element group 735:  members (2) 
      -- CP-element group 735: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/SplitProtocol/Update/$exit
      -- CP-element group 735: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/SplitProtocol/Update/ca
      -- 
    ca_7819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 735_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1859_inst_ack_1, ack => zeropad3D_CP_676_elements(735)); -- 
    -- CP-element group 736:  join  transition  output  bypass 
    -- CP-element group 736: predecessors 
    -- CP-element group 736: 	734 
    -- CP-element group 736: 	735 
    -- CP-element group 736: successors 
    -- CP-element group 736: 	738 
    -- CP-element group 736:  members (5) 
      -- CP-element group 736: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/$exit
      -- CP-element group 736: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/$exit
      -- CP-element group 736: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/$exit
      -- CP-element group 736: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_sources/type_cast_1859/SplitProtocol/$exit
      -- CP-element group 736: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1854/phi_stmt_1854_req
      -- 
    phi_stmt_1854_req_7820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1854_req_7820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(736), ack => phi_stmt_1854_req_1); -- 
    zeropad3D_cp_element_group_736: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_736"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(734) & zeropad3D_CP_676_elements(735);
      gj_zeropad3D_cp_element_group_736 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(736), clk => clk, reset => reset); --
    end block;
    -- CP-element group 737:  transition  output  delay-element  bypass 
    -- CP-element group 737: predecessors 
    -- CP-element group 737: 	284 
    -- CP-element group 737: successors 
    -- CP-element group 737: 	738 
    -- CP-element group 737:  members (4) 
      -- CP-element group 737: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1847/$exit
      -- CP-element group 737: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/$exit
      -- CP-element group 737: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_sources/type_cast_1853_konst_delay_trans
      -- CP-element group 737: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/phi_stmt_1847/phi_stmt_1847_req
      -- 
    phi_stmt_1847_req_7828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1847_req_7828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(737), ack => phi_stmt_1847_req_1); -- 
    -- Element group zeropad3D_CP_676_elements(737) is a control-delay.
    cp_element_737_delay: control_delay_element  generic map(name => " 737_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(284), ack => zeropad3D_CP_676_elements(737), clk => clk, reset =>reset);
    -- CP-element group 738:  join  transition  bypass 
    -- CP-element group 738: predecessors 
    -- CP-element group 738: 	733 
    -- CP-element group 738: 	736 
    -- CP-element group 738: 	737 
    -- CP-element group 738: successors 
    -- CP-element group 738: 	739 
    -- CP-element group 738:  members (1) 
      -- CP-element group 738: 	 branch_block_stmt_223/whilex_xend687_whilex_xbody751_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_738: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_738"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(733) & zeropad3D_CP_676_elements(736) & zeropad3D_CP_676_elements(737);
      gj_zeropad3D_cp_element_group_738 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(738), clk => clk, reset => reset); --
    end block;
    -- CP-element group 739:  merge  fork  transition  place  bypass 
    -- CP-element group 739: predecessors 
    -- CP-element group 739: 	730 
    -- CP-element group 739: 	738 
    -- CP-element group 739: successors 
    -- CP-element group 739: 	740 
    -- CP-element group 739: 	741 
    -- CP-element group 739: 	742 
    -- CP-element group 739:  members (2) 
      -- CP-element group 739: 	 branch_block_stmt_223/merge_stmt_1846_PhiReqMerge
      -- CP-element group 739: 	 branch_block_stmt_223/merge_stmt_1846_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(739) <= OrReduce(zeropad3D_CP_676_elements(730) & zeropad3D_CP_676_elements(738));
    -- CP-element group 740:  transition  input  bypass 
    -- CP-element group 740: predecessors 
    -- CP-element group 740: 	739 
    -- CP-element group 740: successors 
    -- CP-element group 740: 	743 
    -- CP-element group 740:  members (1) 
      -- CP-element group 740: 	 branch_block_stmt_223/merge_stmt_1846_PhiAck/phi_stmt_1847_ack
      -- 
    phi_stmt_1847_ack_7833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 740_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1847_ack_0, ack => zeropad3D_CP_676_elements(740)); -- 
    -- CP-element group 741:  transition  input  bypass 
    -- CP-element group 741: predecessors 
    -- CP-element group 741: 	739 
    -- CP-element group 741: successors 
    -- CP-element group 741: 	743 
    -- CP-element group 741:  members (1) 
      -- CP-element group 741: 	 branch_block_stmt_223/merge_stmt_1846_PhiAck/phi_stmt_1854_ack
      -- 
    phi_stmt_1854_ack_7834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 741_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1854_ack_0, ack => zeropad3D_CP_676_elements(741)); -- 
    -- CP-element group 742:  transition  input  bypass 
    -- CP-element group 742: predecessors 
    -- CP-element group 742: 	739 
    -- CP-element group 742: successors 
    -- CP-element group 742: 	743 
    -- CP-element group 742:  members (1) 
      -- CP-element group 742: 	 branch_block_stmt_223/merge_stmt_1846_PhiAck/phi_stmt_1860_ack
      -- 
    phi_stmt_1860_ack_7835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 742_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1860_ack_0, ack => zeropad3D_CP_676_elements(742)); -- 
    -- CP-element group 743:  join  fork  transition  place  output  bypass 
    -- CP-element group 743: predecessors 
    -- CP-element group 743: 	740 
    -- CP-element group 743: 	741 
    -- CP-element group 743: 	742 
    -- CP-element group 743: successors 
    -- CP-element group 743: 	285 
    -- CP-element group 743: 	286 
    -- CP-element group 743:  members (10) 
      -- CP-element group 743: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896__entry__
      -- CP-element group 743: 	 branch_block_stmt_223/merge_stmt_1846__exit__
      -- CP-element group 743: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/$entry
      -- CP-element group 743: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_sample_start_
      -- CP-element group 743: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_update_start_
      -- CP-element group 743: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_Sample/$entry
      -- CP-element group 743: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_Sample/rr
      -- CP-element group 743: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_Update/$entry
      -- CP-element group 743: 	 branch_block_stmt_223/assign_stmt_1871_to_assign_stmt_1896/type_cast_1870_Update/cr
      -- CP-element group 743: 	 branch_block_stmt_223/merge_stmt_1846_PhiAck/$exit
      -- 
    rr_3633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(743), ack => type_cast_1870_inst_req_0); -- 
    cr_3638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(743), ack => type_cast_1870_inst_req_1); -- 
    zeropad3D_cp_element_group_743: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_743"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(740) & zeropad3D_CP_676_elements(741) & zeropad3D_CP_676_elements(742);
      gj_zeropad3D_cp_element_group_743 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(743), clk => clk, reset => reset); --
    end block;
    -- CP-element group 744:  merge  fork  transition  place  output  bypass 
    -- CP-element group 744: predecessors 
    -- CP-element group 744: 	288 
    -- CP-element group 744: 	292 
    -- CP-element group 744: successors 
    -- CP-element group 744: 	293 
    -- CP-element group 744: 	294 
    -- CP-element group 744: 	295 
    -- CP-element group 744: 	296 
    -- CP-element group 744: 	299 
    -- CP-element group 744: 	301 
    -- CP-element group 744: 	303 
    -- CP-element group 744: 	305 
    -- CP-element group 744:  members (33) 
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996__entry__
      -- CP-element group 744: 	 branch_block_stmt_223/merge_stmt_1940__exit__
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Update/word_access_complete/word_0/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Update/word_access_complete/word_0/cr
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Update/word_access_complete/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_Update/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_sample_start_
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_update_start_
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_Sample/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_Sample/rr
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_Update/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1944_Update/cr
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_sample_start_
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_update_start_
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_Sample/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_Sample/rr
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_Update/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1949_Update/cr
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_update_start_
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_Update/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/type_cast_1983_Update/cr
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_update_start_
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_final_index_sum_regn_update_start
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_final_index_sum_regn_Update/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/array_obj_ref_1989_final_index_sum_regn_Update/req
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_complete/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/addr_of_1990_complete/req
      -- CP-element group 744: 	 branch_block_stmt_223/assign_stmt_1945_to_assign_stmt_1996/ptr_deref_1993_update_start_
      -- CP-element group 744: 	 branch_block_stmt_223/merge_stmt_1940_PhiReqMerge
      -- CP-element group 744: 	 branch_block_stmt_223/merge_stmt_1940_PhiAck/$entry
      -- CP-element group 744: 	 branch_block_stmt_223/merge_stmt_1940_PhiAck/$exit
      -- CP-element group 744: 	 branch_block_stmt_223/merge_stmt_1940_PhiAck/dummy
      -- 
    cr_3834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(744), ack => ptr_deref_1993_store_0_req_1); -- 
    rr_3705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(744), ack => type_cast_1944_inst_req_0); -- 
    cr_3710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(744), ack => type_cast_1944_inst_req_1); -- 
    rr_3719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(744), ack => type_cast_1949_inst_req_0); -- 
    cr_3724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(744), ack => type_cast_1949_inst_req_1); -- 
    cr_3738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(744), ack => type_cast_1983_inst_req_1); -- 
    req_3769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(744), ack => array_obj_ref_1989_index_offset_req_1); -- 
    req_3784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(744), ack => addr_of_1990_final_reg_req_1); -- 
    zeropad3D_CP_676_elements(744) <= OrReduce(zeropad3D_CP_676_elements(288) & zeropad3D_CP_676_elements(292));
    -- CP-element group 745:  merge  fork  transition  place  output  bypass 
    -- CP-element group 745: predecessors 
    -- CP-element group 745: 	306 
    -- CP-element group 745: 	326 
    -- CP-element group 745: successors 
    -- CP-element group 745: 	327 
    -- CP-element group 745: 	328 
    -- CP-element group 745:  members (13) 
      -- CP-element group 745: 	 branch_block_stmt_223/merge_stmt_2105__exit__
      -- CP-element group 745: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123__entry__
      -- CP-element group 745: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_update_start_
      -- CP-element group 745: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_Sample/$entry
      -- CP-element group 745: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_Sample/rr
      -- CP-element group 745: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_Update/$entry
      -- CP-element group 745: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_sample_start_
      -- CP-element group 745: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/$entry
      -- CP-element group 745: 	 branch_block_stmt_223/assign_stmt_2110_to_assign_stmt_2123/type_cast_2109_Update/cr
      -- CP-element group 745: 	 branch_block_stmt_223/merge_stmt_2105_PhiReqMerge
      -- CP-element group 745: 	 branch_block_stmt_223/merge_stmt_2105_PhiAck/$entry
      -- CP-element group 745: 	 branch_block_stmt_223/merge_stmt_2105_PhiAck/$exit
      -- CP-element group 745: 	 branch_block_stmt_223/merge_stmt_2105_PhiAck/dummy
      -- 
    rr_4083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(745), ack => type_cast_2109_inst_req_0); -- 
    cr_4088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(745), ack => type_cast_2109_inst_req_1); -- 
    zeropad3D_CP_676_elements(745) <= OrReduce(zeropad3D_CP_676_elements(306) & zeropad3D_CP_676_elements(326));
    -- CP-element group 746:  transition  output  delay-element  bypass 
    -- CP-element group 746: predecessors 
    -- CP-element group 746: 	338 
    -- CP-element group 746: successors 
    -- CP-element group 746: 	753 
    -- CP-element group 746:  members (4) 
      -- CP-element group 746: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2187/$exit
      -- CP-element group 746: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/$exit
      -- CP-element group 746: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2191_konst_delay_trans
      -- CP-element group 746: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_req
      -- 
    phi_stmt_2187_req_7916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2187_req_7916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(746), ack => phi_stmt_2187_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(746) is a control-delay.
    cp_element_746_delay: control_delay_element  generic map(name => " 746_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(338), ack => zeropad3D_CP_676_elements(746), clk => clk, reset =>reset);
    -- CP-element group 747:  transition  input  bypass 
    -- CP-element group 747: predecessors 
    -- CP-element group 747: 	338 
    -- CP-element group 747: successors 
    -- CP-element group 747: 	749 
    -- CP-element group 747:  members (2) 
      -- CP-element group 747: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/$exit
      -- CP-element group 747: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/ra
      -- 
    ra_7933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 747_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_0, ack => zeropad3D_CP_676_elements(747)); -- 
    -- CP-element group 748:  transition  input  bypass 
    -- CP-element group 748: predecessors 
    -- CP-element group 748: 	338 
    -- CP-element group 748: successors 
    -- CP-element group 748: 	749 
    -- CP-element group 748:  members (2) 
      -- CP-element group 748: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/$exit
      -- CP-element group 748: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/ca
      -- 
    ca_7938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 748_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_1, ack => zeropad3D_CP_676_elements(748)); -- 
    -- CP-element group 749:  join  transition  output  bypass 
    -- CP-element group 749: predecessors 
    -- CP-element group 749: 	747 
    -- CP-element group 749: 	748 
    -- CP-element group 749: successors 
    -- CP-element group 749: 	753 
    -- CP-element group 749:  members (5) 
      -- CP-element group 749: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/$exit
      -- CP-element group 749: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$exit
      -- CP-element group 749: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/$exit
      -- CP-element group 749: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/$exit
      -- CP-element group 749: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_req
      -- 
    phi_stmt_2194_req_7939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2194_req_7939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(749), ack => phi_stmt_2194_req_1); -- 
    zeropad3D_cp_element_group_749: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_749"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(747) & zeropad3D_CP_676_elements(748);
      gj_zeropad3D_cp_element_group_749 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(749), clk => clk, reset => reset); --
    end block;
    -- CP-element group 750:  transition  input  bypass 
    -- CP-element group 750: predecessors 
    -- CP-element group 750: 	338 
    -- CP-element group 750: successors 
    -- CP-element group 750: 	752 
    -- CP-element group 750:  members (2) 
      -- CP-element group 750: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/SplitProtocol/Sample/$exit
      -- CP-element group 750: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/SplitProtocol/Sample/ra
      -- 
    ra_7956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 750_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2203_inst_ack_0, ack => zeropad3D_CP_676_elements(750)); -- 
    -- CP-element group 751:  transition  input  bypass 
    -- CP-element group 751: predecessors 
    -- CP-element group 751: 	338 
    -- CP-element group 751: successors 
    -- CP-element group 751: 	752 
    -- CP-element group 751:  members (2) 
      -- CP-element group 751: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/SplitProtocol/Update/$exit
      -- CP-element group 751: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/SplitProtocol/Update/ca
      -- 
    ca_7961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 751_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2203_inst_ack_1, ack => zeropad3D_CP_676_elements(751)); -- 
    -- CP-element group 752:  join  transition  output  bypass 
    -- CP-element group 752: predecessors 
    -- CP-element group 752: 	750 
    -- CP-element group 752: 	751 
    -- CP-element group 752: successors 
    -- CP-element group 752: 	753 
    -- CP-element group 752:  members (5) 
      -- CP-element group 752: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/$exit
      -- CP-element group 752: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/$exit
      -- CP-element group 752: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/$exit
      -- CP-element group 752: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2203/SplitProtocol/$exit
      -- CP-element group 752: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_req
      -- 
    phi_stmt_2200_req_7962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2200_req_7962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(752), ack => phi_stmt_2200_req_0); -- 
    zeropad3D_cp_element_group_752: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_752"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(750) & zeropad3D_CP_676_elements(751);
      gj_zeropad3D_cp_element_group_752 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(752), clk => clk, reset => reset); --
    end block;
    -- CP-element group 753:  join  transition  bypass 
    -- CP-element group 753: predecessors 
    -- CP-element group 753: 	746 
    -- CP-element group 753: 	749 
    -- CP-element group 753: 	752 
    -- CP-element group 753: successors 
    -- CP-element group 753: 	764 
    -- CP-element group 753:  members (1) 
      -- CP-element group 753: 	 branch_block_stmt_223/ifx_xelse870_ifx_xend906_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_753: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_753"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(746) & zeropad3D_CP_676_elements(749) & zeropad3D_CP_676_elements(752);
      gj_zeropad3D_cp_element_group_753 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(753), clk => clk, reset => reset); --
    end block;
    -- CP-element group 754:  transition  input  bypass 
    -- CP-element group 754: predecessors 
    -- CP-element group 754: 	329 
    -- CP-element group 754: successors 
    -- CP-element group 754: 	756 
    -- CP-element group 754:  members (2) 
      -- CP-element group 754: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/SplitProtocol/Sample/$exit
      -- CP-element group 754: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/SplitProtocol/Sample/ra
      -- 
    ra_7982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 754_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_0, ack => zeropad3D_CP_676_elements(754)); -- 
    -- CP-element group 755:  transition  input  bypass 
    -- CP-element group 755: predecessors 
    -- CP-element group 755: 	329 
    -- CP-element group 755: successors 
    -- CP-element group 755: 	756 
    -- CP-element group 755:  members (2) 
      -- CP-element group 755: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/SplitProtocol/Update/$exit
      -- CP-element group 755: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/SplitProtocol/Update/ca
      -- 
    ca_7987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 755_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_1, ack => zeropad3D_CP_676_elements(755)); -- 
    -- CP-element group 756:  join  transition  output  bypass 
    -- CP-element group 756: predecessors 
    -- CP-element group 756: 	754 
    -- CP-element group 756: 	755 
    -- CP-element group 756: successors 
    -- CP-element group 756: 	763 
    -- CP-element group 756:  members (5) 
      -- CP-element group 756: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/$exit
      -- CP-element group 756: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/$exit
      -- CP-element group 756: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/$exit
      -- CP-element group 756: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193/SplitProtocol/$exit
      -- CP-element group 756: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2187/phi_stmt_2187_req
      -- 
    phi_stmt_2187_req_7988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2187_req_7988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(756), ack => phi_stmt_2187_req_1); -- 
    zeropad3D_cp_element_group_756: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_756"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(754) & zeropad3D_CP_676_elements(755);
      gj_zeropad3D_cp_element_group_756 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(756), clk => clk, reset => reset); --
    end block;
    -- CP-element group 757:  transition  input  bypass 
    -- CP-element group 757: predecessors 
    -- CP-element group 757: 	329 
    -- CP-element group 757: successors 
    -- CP-element group 757: 	759 
    -- CP-element group 757:  members (2) 
      -- CP-element group 757: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/$exit
      -- CP-element group 757: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/ra
      -- 
    ra_8005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 757_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2197_inst_ack_0, ack => zeropad3D_CP_676_elements(757)); -- 
    -- CP-element group 758:  transition  input  bypass 
    -- CP-element group 758: predecessors 
    -- CP-element group 758: 	329 
    -- CP-element group 758: successors 
    -- CP-element group 758: 	759 
    -- CP-element group 758:  members (2) 
      -- CP-element group 758: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/$exit
      -- CP-element group 758: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/ca
      -- 
    ca_8010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 758_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2197_inst_ack_1, ack => zeropad3D_CP_676_elements(758)); -- 
    -- CP-element group 759:  join  transition  output  bypass 
    -- CP-element group 759: predecessors 
    -- CP-element group 759: 	757 
    -- CP-element group 759: 	758 
    -- CP-element group 759: successors 
    -- CP-element group 759: 	763 
    -- CP-element group 759:  members (5) 
      -- CP-element group 759: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/$exit
      -- CP-element group 759: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$exit
      -- CP-element group 759: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/$exit
      -- CP-element group 759: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/$exit
      -- CP-element group 759: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2194/phi_stmt_2194_req
      -- 
    phi_stmt_2194_req_8011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2194_req_8011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(759), ack => phi_stmt_2194_req_0); -- 
    zeropad3D_cp_element_group_759: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_759"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(757) & zeropad3D_CP_676_elements(758);
      gj_zeropad3D_cp_element_group_759 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(759), clk => clk, reset => reset); --
    end block;
    -- CP-element group 760:  transition  input  bypass 
    -- CP-element group 760: predecessors 
    -- CP-element group 760: 	329 
    -- CP-element group 760: successors 
    -- CP-element group 760: 	762 
    -- CP-element group 760:  members (2) 
      -- CP-element group 760: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/SplitProtocol/Sample/$exit
      -- CP-element group 760: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/SplitProtocol/Sample/ra
      -- 
    ra_8028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 760_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2205_inst_ack_0, ack => zeropad3D_CP_676_elements(760)); -- 
    -- CP-element group 761:  transition  input  bypass 
    -- CP-element group 761: predecessors 
    -- CP-element group 761: 	329 
    -- CP-element group 761: successors 
    -- CP-element group 761: 	762 
    -- CP-element group 761:  members (2) 
      -- CP-element group 761: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/SplitProtocol/Update/$exit
      -- CP-element group 761: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/SplitProtocol/Update/ca
      -- 
    ca_8033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 761_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2205_inst_ack_1, ack => zeropad3D_CP_676_elements(761)); -- 
    -- CP-element group 762:  join  transition  output  bypass 
    -- CP-element group 762: predecessors 
    -- CP-element group 762: 	760 
    -- CP-element group 762: 	761 
    -- CP-element group 762: successors 
    -- CP-element group 762: 	763 
    -- CP-element group 762:  members (5) 
      -- CP-element group 762: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/$exit
      -- CP-element group 762: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/$exit
      -- CP-element group 762: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/$exit
      -- CP-element group 762: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_sources/type_cast_2205/SplitProtocol/$exit
      -- CP-element group 762: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/phi_stmt_2200/phi_stmt_2200_req
      -- 
    phi_stmt_2200_req_8034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2200_req_8034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(762), ack => phi_stmt_2200_req_1); -- 
    zeropad3D_cp_element_group_762: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_762"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(760) & zeropad3D_CP_676_elements(761);
      gj_zeropad3D_cp_element_group_762 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(762), clk => clk, reset => reset); --
    end block;
    -- CP-element group 763:  join  transition  bypass 
    -- CP-element group 763: predecessors 
    -- CP-element group 763: 	756 
    -- CP-element group 763: 	759 
    -- CP-element group 763: 	762 
    -- CP-element group 763: successors 
    -- CP-element group 763: 	764 
    -- CP-element group 763:  members (1) 
      -- CP-element group 763: 	 branch_block_stmt_223/ifx_xthen865_ifx_xend906_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_763: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_763"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(756) & zeropad3D_CP_676_elements(759) & zeropad3D_CP_676_elements(762);
      gj_zeropad3D_cp_element_group_763 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(763), clk => clk, reset => reset); --
    end block;
    -- CP-element group 764:  merge  fork  transition  place  bypass 
    -- CP-element group 764: predecessors 
    -- CP-element group 764: 	753 
    -- CP-element group 764: 	763 
    -- CP-element group 764: successors 
    -- CP-element group 764: 	765 
    -- CP-element group 764: 	766 
    -- CP-element group 764: 	767 
    -- CP-element group 764:  members (2) 
      -- CP-element group 764: 	 branch_block_stmt_223/merge_stmt_2186_PhiReqMerge
      -- CP-element group 764: 	 branch_block_stmt_223/merge_stmt_2186_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(764) <= OrReduce(zeropad3D_CP_676_elements(753) & zeropad3D_CP_676_elements(763));
    -- CP-element group 765:  transition  input  bypass 
    -- CP-element group 765: predecessors 
    -- CP-element group 765: 	764 
    -- CP-element group 765: successors 
    -- CP-element group 765: 	768 
    -- CP-element group 765:  members (1) 
      -- CP-element group 765: 	 branch_block_stmt_223/merge_stmt_2186_PhiAck/phi_stmt_2187_ack
      -- 
    phi_stmt_2187_ack_8039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 765_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2187_ack_0, ack => zeropad3D_CP_676_elements(765)); -- 
    -- CP-element group 766:  transition  input  bypass 
    -- CP-element group 766: predecessors 
    -- CP-element group 766: 	764 
    -- CP-element group 766: successors 
    -- CP-element group 766: 	768 
    -- CP-element group 766:  members (1) 
      -- CP-element group 766: 	 branch_block_stmt_223/merge_stmt_2186_PhiAck/phi_stmt_2194_ack
      -- 
    phi_stmt_2194_ack_8040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 766_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2194_ack_0, ack => zeropad3D_CP_676_elements(766)); -- 
    -- CP-element group 767:  transition  input  bypass 
    -- CP-element group 767: predecessors 
    -- CP-element group 767: 	764 
    -- CP-element group 767: successors 
    -- CP-element group 767: 	768 
    -- CP-element group 767:  members (1) 
      -- CP-element group 767: 	 branch_block_stmt_223/merge_stmt_2186_PhiAck/phi_stmt_2200_ack
      -- 
    phi_stmt_2200_ack_8041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 767_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2200_ack_0, ack => zeropad3D_CP_676_elements(767)); -- 
    -- CP-element group 768:  join  transition  bypass 
    -- CP-element group 768: predecessors 
    -- CP-element group 768: 	765 
    -- CP-element group 768: 	766 
    -- CP-element group 768: 	767 
    -- CP-element group 768: successors 
    -- CP-element group 768: 	4 
    -- CP-element group 768:  members (1) 
      -- CP-element group 768: 	 branch_block_stmt_223/merge_stmt_2186_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_768: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_768"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(765) & zeropad3D_CP_676_elements(766) & zeropad3D_CP_676_elements(767);
      gj_zeropad3D_cp_element_group_768 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(768), clk => clk, reset => reset); --
    end block;
    -- CP-element group 769:  transition  input  bypass 
    -- CP-element group 769: predecessors 
    -- CP-element group 769: 	5 
    -- CP-element group 769: successors 
    -- CP-element group 769: 	771 
    -- CP-element group 769:  members (2) 
      -- CP-element group 769: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/SplitProtocol/Sample/$exit
      -- CP-element group 769: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/SplitProtocol/Sample/ra
      -- 
    ra_8069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 769_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2268_inst_ack_0, ack => zeropad3D_CP_676_elements(769)); -- 
    -- CP-element group 770:  transition  input  bypass 
    -- CP-element group 770: predecessors 
    -- CP-element group 770: 	5 
    -- CP-element group 770: successors 
    -- CP-element group 770: 	771 
    -- CP-element group 770:  members (2) 
      -- CP-element group 770: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/SplitProtocol/Update/$exit
      -- CP-element group 770: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/SplitProtocol/Update/ca
      -- 
    ca_8074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 770_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2268_inst_ack_1, ack => zeropad3D_CP_676_elements(770)); -- 
    -- CP-element group 771:  join  transition  output  bypass 
    -- CP-element group 771: predecessors 
    -- CP-element group 771: 	769 
    -- CP-element group 771: 	770 
    -- CP-element group 771: successors 
    -- CP-element group 771: 	778 
    -- CP-element group 771:  members (5) 
      -- CP-element group 771: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/$exit
      -- CP-element group 771: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/$exit
      -- CP-element group 771: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/$exit
      -- CP-element group 771: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2268/SplitProtocol/$exit
      -- CP-element group 771: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_req
      -- 
    phi_stmt_2262_req_8075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2262_req_8075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(771), ack => phi_stmt_2262_req_1); -- 
    zeropad3D_cp_element_group_771: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_771"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(769) & zeropad3D_CP_676_elements(770);
      gj_zeropad3D_cp_element_group_771 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(771), clk => clk, reset => reset); --
    end block;
    -- CP-element group 772:  transition  input  bypass 
    -- CP-element group 772: predecessors 
    -- CP-element group 772: 	5 
    -- CP-element group 772: successors 
    -- CP-element group 772: 	774 
    -- CP-element group 772:  members (2) 
      -- CP-element group 772: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/SplitProtocol/Sample/$exit
      -- CP-element group 772: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/SplitProtocol/Sample/ra
      -- 
    ra_8092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 772_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2274_inst_ack_0, ack => zeropad3D_CP_676_elements(772)); -- 
    -- CP-element group 773:  transition  input  bypass 
    -- CP-element group 773: predecessors 
    -- CP-element group 773: 	5 
    -- CP-element group 773: successors 
    -- CP-element group 773: 	774 
    -- CP-element group 773:  members (2) 
      -- CP-element group 773: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/SplitProtocol/Update/$exit
      -- CP-element group 773: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/SplitProtocol/Update/ca
      -- 
    ca_8097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 773_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2274_inst_ack_1, ack => zeropad3D_CP_676_elements(773)); -- 
    -- CP-element group 774:  join  transition  output  bypass 
    -- CP-element group 774: predecessors 
    -- CP-element group 774: 	772 
    -- CP-element group 774: 	773 
    -- CP-element group 774: successors 
    -- CP-element group 774: 	778 
    -- CP-element group 774:  members (5) 
      -- CP-element group 774: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/$exit
      -- CP-element group 774: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/$exit
      -- CP-element group 774: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/$exit
      -- CP-element group 774: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2274/SplitProtocol/$exit
      -- CP-element group 774: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_req
      -- 
    phi_stmt_2269_req_8098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2269_req_8098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(774), ack => phi_stmt_2269_req_1); -- 
    zeropad3D_cp_element_group_774: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_774"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(772) & zeropad3D_CP_676_elements(773);
      gj_zeropad3D_cp_element_group_774 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(774), clk => clk, reset => reset); --
    end block;
    -- CP-element group 775:  transition  input  bypass 
    -- CP-element group 775: predecessors 
    -- CP-element group 775: 	5 
    -- CP-element group 775: successors 
    -- CP-element group 775: 	777 
    -- CP-element group 775:  members (2) 
      -- CP-element group 775: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/SplitProtocol/Sample/$exit
      -- CP-element group 775: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/SplitProtocol/Sample/ra
      -- 
    ra_8115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 775_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2281_inst_ack_0, ack => zeropad3D_CP_676_elements(775)); -- 
    -- CP-element group 776:  transition  input  bypass 
    -- CP-element group 776: predecessors 
    -- CP-element group 776: 	5 
    -- CP-element group 776: successors 
    -- CP-element group 776: 	777 
    -- CP-element group 776:  members (2) 
      -- CP-element group 776: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/SplitProtocol/Update/$exit
      -- CP-element group 776: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/SplitProtocol/Update/ca
      -- 
    ca_8120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 776_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2281_inst_ack_1, ack => zeropad3D_CP_676_elements(776)); -- 
    -- CP-element group 777:  join  transition  output  bypass 
    -- CP-element group 777: predecessors 
    -- CP-element group 777: 	775 
    -- CP-element group 777: 	776 
    -- CP-element group 777: successors 
    -- CP-element group 777: 	778 
    -- CP-element group 777:  members (5) 
      -- CP-element group 777: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/$exit
      -- CP-element group 777: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/$exit
      -- CP-element group 777: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/$exit
      -- CP-element group 777: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2281/SplitProtocol/$exit
      -- CP-element group 777: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_req
      -- 
    phi_stmt_2275_req_8121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2275_req_8121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(777), ack => phi_stmt_2275_req_1); -- 
    zeropad3D_cp_element_group_777: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_777"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(775) & zeropad3D_CP_676_elements(776);
      gj_zeropad3D_cp_element_group_777 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(777), clk => clk, reset => reset); --
    end block;
    -- CP-element group 778:  join  transition  bypass 
    -- CP-element group 778: predecessors 
    -- CP-element group 778: 	771 
    -- CP-element group 778: 	774 
    -- CP-element group 778: 	777 
    -- CP-element group 778: successors 
    -- CP-element group 778: 	785 
    -- CP-element group 778:  members (1) 
      -- CP-element group 778: 	 branch_block_stmt_223/ifx_xend1126_whilex_xbody967_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_778: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_778"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(771) & zeropad3D_CP_676_elements(774) & zeropad3D_CP_676_elements(777);
      gj_zeropad3D_cp_element_group_778 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(778), clk => clk, reset => reset); --
    end block;
    -- CP-element group 779:  transition  output  delay-element  bypass 
    -- CP-element group 779: predecessors 
    -- CP-element group 779: 	342 
    -- CP-element group 779: successors 
    -- CP-element group 779: 	784 
    -- CP-element group 779:  members (4) 
      -- CP-element group 779: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2262/$exit
      -- CP-element group 779: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/$exit
      -- CP-element group 779: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_sources/type_cast_2266_konst_delay_trans
      -- CP-element group 779: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2262/phi_stmt_2262_req
      -- 
    phi_stmt_2262_req_8132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2262_req_8132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(779), ack => phi_stmt_2262_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(779) is a control-delay.
    cp_element_779_delay: control_delay_element  generic map(name => " 779_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(342), ack => zeropad3D_CP_676_elements(779), clk => clk, reset =>reset);
    -- CP-element group 780:  transition  input  bypass 
    -- CP-element group 780: predecessors 
    -- CP-element group 780: 	342 
    -- CP-element group 780: successors 
    -- CP-element group 780: 	782 
    -- CP-element group 780:  members (2) 
      -- CP-element group 780: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Sample/$exit
      -- CP-element group 780: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Sample/ra
      -- 
    ra_8149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 780_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2272_inst_ack_0, ack => zeropad3D_CP_676_elements(780)); -- 
    -- CP-element group 781:  transition  input  bypass 
    -- CP-element group 781: predecessors 
    -- CP-element group 781: 	342 
    -- CP-element group 781: successors 
    -- CP-element group 781: 	782 
    -- CP-element group 781:  members (2) 
      -- CP-element group 781: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Update/$exit
      -- CP-element group 781: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/Update/ca
      -- 
    ca_8154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 781_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2272_inst_ack_1, ack => zeropad3D_CP_676_elements(781)); -- 
    -- CP-element group 782:  join  transition  output  bypass 
    -- CP-element group 782: predecessors 
    -- CP-element group 782: 	780 
    -- CP-element group 782: 	781 
    -- CP-element group 782: successors 
    -- CP-element group 782: 	784 
    -- CP-element group 782:  members (5) 
      -- CP-element group 782: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/$exit
      -- CP-element group 782: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/$exit
      -- CP-element group 782: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/$exit
      -- CP-element group 782: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_sources/type_cast_2272/SplitProtocol/$exit
      -- CP-element group 782: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2269/phi_stmt_2269_req
      -- 
    phi_stmt_2269_req_8155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2269_req_8155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(782), ack => phi_stmt_2269_req_0); -- 
    zeropad3D_cp_element_group_782: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_782"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(780) & zeropad3D_CP_676_elements(781);
      gj_zeropad3D_cp_element_group_782 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(782), clk => clk, reset => reset); --
    end block;
    -- CP-element group 783:  transition  output  delay-element  bypass 
    -- CP-element group 783: predecessors 
    -- CP-element group 783: 	342 
    -- CP-element group 783: successors 
    -- CP-element group 783: 	784 
    -- CP-element group 783:  members (4) 
      -- CP-element group 783: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2275/$exit
      -- CP-element group 783: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/$exit
      -- CP-element group 783: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_sources/type_cast_2279_konst_delay_trans
      -- CP-element group 783: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/phi_stmt_2275/phi_stmt_2275_req
      -- 
    phi_stmt_2275_req_8163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2275_req_8163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(783), ack => phi_stmt_2275_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(783) is a control-delay.
    cp_element_783_delay: control_delay_element  generic map(name => " 783_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(342), ack => zeropad3D_CP_676_elements(783), clk => clk, reset =>reset);
    -- CP-element group 784:  join  transition  bypass 
    -- CP-element group 784: predecessors 
    -- CP-element group 784: 	779 
    -- CP-element group 784: 	782 
    -- CP-element group 784: 	783 
    -- CP-element group 784: successors 
    -- CP-element group 784: 	785 
    -- CP-element group 784:  members (1) 
      -- CP-element group 784: 	 branch_block_stmt_223/whilex_xend907_whilex_xbody967_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_784: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_784"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(779) & zeropad3D_CP_676_elements(782) & zeropad3D_CP_676_elements(783);
      gj_zeropad3D_cp_element_group_784 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(784), clk => clk, reset => reset); --
    end block;
    -- CP-element group 785:  merge  fork  transition  place  bypass 
    -- CP-element group 785: predecessors 
    -- CP-element group 785: 	778 
    -- CP-element group 785: 	784 
    -- CP-element group 785: successors 
    -- CP-element group 785: 	786 
    -- CP-element group 785: 	787 
    -- CP-element group 785: 	788 
    -- CP-element group 785:  members (2) 
      -- CP-element group 785: 	 branch_block_stmt_223/merge_stmt_2261_PhiReqMerge
      -- CP-element group 785: 	 branch_block_stmt_223/merge_stmt_2261_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(785) <= OrReduce(zeropad3D_CP_676_elements(778) & zeropad3D_CP_676_elements(784));
    -- CP-element group 786:  transition  input  bypass 
    -- CP-element group 786: predecessors 
    -- CP-element group 786: 	785 
    -- CP-element group 786: successors 
    -- CP-element group 786: 	789 
    -- CP-element group 786:  members (1) 
      -- CP-element group 786: 	 branch_block_stmt_223/merge_stmt_2261_PhiAck/phi_stmt_2262_ack
      -- 
    phi_stmt_2262_ack_8168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 786_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2262_ack_0, ack => zeropad3D_CP_676_elements(786)); -- 
    -- CP-element group 787:  transition  input  bypass 
    -- CP-element group 787: predecessors 
    -- CP-element group 787: 	785 
    -- CP-element group 787: successors 
    -- CP-element group 787: 	789 
    -- CP-element group 787:  members (1) 
      -- CP-element group 787: 	 branch_block_stmt_223/merge_stmt_2261_PhiAck/phi_stmt_2269_ack
      -- 
    phi_stmt_2269_ack_8169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 787_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2269_ack_0, ack => zeropad3D_CP_676_elements(787)); -- 
    -- CP-element group 788:  transition  input  bypass 
    -- CP-element group 788: predecessors 
    -- CP-element group 788: 	785 
    -- CP-element group 788: successors 
    -- CP-element group 788: 	789 
    -- CP-element group 788:  members (1) 
      -- CP-element group 788: 	 branch_block_stmt_223/merge_stmt_2261_PhiAck/phi_stmt_2275_ack
      -- 
    phi_stmt_2275_ack_8170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 788_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2275_ack_0, ack => zeropad3D_CP_676_elements(788)); -- 
    -- CP-element group 789:  join  fork  transition  place  output  bypass 
    -- CP-element group 789: predecessors 
    -- CP-element group 789: 	786 
    -- CP-element group 789: 	787 
    -- CP-element group 789: 	788 
    -- CP-element group 789: successors 
    -- CP-element group 789: 	343 
    -- CP-element group 789: 	344 
    -- CP-element group 789:  members (10) 
      -- CP-element group 789: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312__entry__
      -- CP-element group 789: 	 branch_block_stmt_223/merge_stmt_2261__exit__
      -- CP-element group 789: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/$entry
      -- CP-element group 789: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_sample_start_
      -- CP-element group 789: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_update_start_
      -- CP-element group 789: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_Sample/$entry
      -- CP-element group 789: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_Sample/rr
      -- CP-element group 789: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_Update/$entry
      -- CP-element group 789: 	 branch_block_stmt_223/assign_stmt_2287_to_assign_stmt_2312/type_cast_2286_Update/cr
      -- CP-element group 789: 	 branch_block_stmt_223/merge_stmt_2261_PhiAck/$exit
      -- 
    rr_4236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(789), ack => type_cast_2286_inst_req_0); -- 
    cr_4241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(789), ack => type_cast_2286_inst_req_1); -- 
    zeropad3D_cp_element_group_789: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_789"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(786) & zeropad3D_CP_676_elements(787) & zeropad3D_CP_676_elements(788);
      gj_zeropad3D_cp_element_group_789 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(789), clk => clk, reset => reset); --
    end block;
    -- CP-element group 790:  merge  fork  transition  place  output  bypass 
    -- CP-element group 790: predecessors 
    -- CP-element group 790: 	346 
    -- CP-element group 790: 	350 
    -- CP-element group 790: successors 
    -- CP-element group 790: 	351 
    -- CP-element group 790: 	352 
    -- CP-element group 790: 	353 
    -- CP-element group 790: 	354 
    -- CP-element group 790: 	357 
    -- CP-element group 790: 	359 
    -- CP-element group 790: 	361 
    -- CP-element group 790: 	363 
    -- CP-element group 790:  members (33) 
      -- CP-element group 790: 	 branch_block_stmt_223/merge_stmt_2356__exit__
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412__entry__
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_sample_start_
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_update_start_
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_Sample/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_Sample/rr
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_Update/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2360_Update/cr
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_sample_start_
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_update_start_
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_Sample/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_Sample/rr
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_Update/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2365_Update/cr
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_update_start_
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_Update/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/type_cast_2399_Update/cr
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_update_start_
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_final_index_sum_regn_update_start
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_final_index_sum_regn_Update/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/array_obj_ref_2405_final_index_sum_regn_Update/req
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_complete/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/addr_of_2406_complete/req
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_update_start_
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Update/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Update/word_access_complete/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Update/word_access_complete/word_0/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/assign_stmt_2361_to_assign_stmt_2412/ptr_deref_2409_Update/word_access_complete/word_0/cr
      -- CP-element group 790: 	 branch_block_stmt_223/merge_stmt_2356_PhiReqMerge
      -- CP-element group 790: 	 branch_block_stmt_223/merge_stmt_2356_PhiAck/$entry
      -- CP-element group 790: 	 branch_block_stmt_223/merge_stmt_2356_PhiAck/$exit
      -- CP-element group 790: 	 branch_block_stmt_223/merge_stmt_2356_PhiAck/dummy
      -- 
    rr_4308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(790), ack => type_cast_2360_inst_req_0); -- 
    cr_4313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(790), ack => type_cast_2360_inst_req_1); -- 
    rr_4322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(790), ack => type_cast_2365_inst_req_0); -- 
    cr_4327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(790), ack => type_cast_2365_inst_req_1); -- 
    cr_4341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(790), ack => type_cast_2399_inst_req_1); -- 
    req_4372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(790), ack => array_obj_ref_2405_index_offset_req_1); -- 
    req_4387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(790), ack => addr_of_2406_final_reg_req_1); -- 
    cr_4437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(790), ack => ptr_deref_2409_store_0_req_1); -- 
    zeropad3D_CP_676_elements(790) <= OrReduce(zeropad3D_CP_676_elements(346) & zeropad3D_CP_676_elements(350));
    -- CP-element group 791:  merge  fork  transition  place  output  bypass 
    -- CP-element group 791: predecessors 
    -- CP-element group 791: 	364 
    -- CP-element group 791: 	384 
    -- CP-element group 791: successors 
    -- CP-element group 791: 	385 
    -- CP-element group 791: 	386 
    -- CP-element group 791:  members (13) 
      -- CP-element group 791: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539__entry__
      -- CP-element group 791: 	 branch_block_stmt_223/merge_stmt_2521__exit__
      -- CP-element group 791: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/$entry
      -- CP-element group 791: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_sample_start_
      -- CP-element group 791: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_update_start_
      -- CP-element group 791: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_Sample/$entry
      -- CP-element group 791: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_Sample/rr
      -- CP-element group 791: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_Update/$entry
      -- CP-element group 791: 	 branch_block_stmt_223/assign_stmt_2526_to_assign_stmt_2539/type_cast_2525_Update/cr
      -- CP-element group 791: 	 branch_block_stmt_223/merge_stmt_2521_PhiReqMerge
      -- CP-element group 791: 	 branch_block_stmt_223/merge_stmt_2521_PhiAck/$entry
      -- CP-element group 791: 	 branch_block_stmt_223/merge_stmt_2521_PhiAck/$exit
      -- CP-element group 791: 	 branch_block_stmt_223/merge_stmt_2521_PhiAck/dummy
      -- 
    rr_4686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(791), ack => type_cast_2525_inst_req_0); -- 
    cr_4691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(791), ack => type_cast_2525_inst_req_1); -- 
    zeropad3D_CP_676_elements(791) <= OrReduce(zeropad3D_CP_676_elements(364) & zeropad3D_CP_676_elements(384));
    -- CP-element group 792:  transition  output  delay-element  bypass 
    -- CP-element group 792: predecessors 
    -- CP-element group 792: 	396 
    -- CP-element group 792: successors 
    -- CP-element group 792: 	799 
    -- CP-element group 792:  members (4) 
      -- CP-element group 792: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2604/$exit
      -- CP-element group 792: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/$exit
      -- CP-element group 792: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2610_konst_delay_trans
      -- CP-element group 792: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_req
      -- 
    phi_stmt_2604_req_8251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2604_req_8251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(792), ack => phi_stmt_2604_req_1); -- 
    -- Element group zeropad3D_CP_676_elements(792) is a control-delay.
    cp_element_792_delay: control_delay_element  generic map(name => " 792_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(396), ack => zeropad3D_CP_676_elements(792), clk => clk, reset =>reset);
    -- CP-element group 793:  transition  input  bypass 
    -- CP-element group 793: predecessors 
    -- CP-element group 793: 	396 
    -- CP-element group 793: successors 
    -- CP-element group 793: 	795 
    -- CP-element group 793:  members (2) 
      -- CP-element group 793: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/SplitProtocol/Sample/$exit
      -- CP-element group 793: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/SplitProtocol/Sample/ra
      -- 
    ra_8268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 793_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2616_inst_ack_0, ack => zeropad3D_CP_676_elements(793)); -- 
    -- CP-element group 794:  transition  input  bypass 
    -- CP-element group 794: predecessors 
    -- CP-element group 794: 	396 
    -- CP-element group 794: successors 
    -- CP-element group 794: 	795 
    -- CP-element group 794:  members (2) 
      -- CP-element group 794: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/SplitProtocol/Update/$exit
      -- CP-element group 794: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/SplitProtocol/Update/ca
      -- 
    ca_8273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 794_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2616_inst_ack_1, ack => zeropad3D_CP_676_elements(794)); -- 
    -- CP-element group 795:  join  transition  output  bypass 
    -- CP-element group 795: predecessors 
    -- CP-element group 795: 	793 
    -- CP-element group 795: 	794 
    -- CP-element group 795: successors 
    -- CP-element group 795: 	799 
    -- CP-element group 795:  members (5) 
      -- CP-element group 795: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/$exit
      -- CP-element group 795: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/$exit
      -- CP-element group 795: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/$exit
      -- CP-element group 795: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2616/SplitProtocol/$exit
      -- CP-element group 795: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_req
      -- 
    phi_stmt_2611_req_8274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2611_req_8274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(795), ack => phi_stmt_2611_req_1); -- 
    zeropad3D_cp_element_group_795: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_795"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(793) & zeropad3D_CP_676_elements(794);
      gj_zeropad3D_cp_element_group_795 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(795), clk => clk, reset => reset); --
    end block;
    -- CP-element group 796:  transition  input  bypass 
    -- CP-element group 796: predecessors 
    -- CP-element group 796: 	396 
    -- CP-element group 796: successors 
    -- CP-element group 796: 	798 
    -- CP-element group 796:  members (2) 
      -- CP-element group 796: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/SplitProtocol/Sample/$exit
      -- CP-element group 796: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/SplitProtocol/Sample/ra
      -- 
    ra_8291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 796_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2622_inst_ack_0, ack => zeropad3D_CP_676_elements(796)); -- 
    -- CP-element group 797:  transition  input  bypass 
    -- CP-element group 797: predecessors 
    -- CP-element group 797: 	396 
    -- CP-element group 797: successors 
    -- CP-element group 797: 	798 
    -- CP-element group 797:  members (2) 
      -- CP-element group 797: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/SplitProtocol/Update/$exit
      -- CP-element group 797: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/SplitProtocol/Update/ca
      -- 
    ca_8296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 797_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2622_inst_ack_1, ack => zeropad3D_CP_676_elements(797)); -- 
    -- CP-element group 798:  join  transition  output  bypass 
    -- CP-element group 798: predecessors 
    -- CP-element group 798: 	796 
    -- CP-element group 798: 	797 
    -- CP-element group 798: successors 
    -- CP-element group 798: 	799 
    -- CP-element group 798:  members (5) 
      -- CP-element group 798: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/$exit
      -- CP-element group 798: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/$exit
      -- CP-element group 798: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/$exit
      -- CP-element group 798: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2622/SplitProtocol/$exit
      -- CP-element group 798: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_req
      -- 
    phi_stmt_2617_req_8297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2617_req_8297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(798), ack => phi_stmt_2617_req_1); -- 
    zeropad3D_cp_element_group_798: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_798"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(796) & zeropad3D_CP_676_elements(797);
      gj_zeropad3D_cp_element_group_798 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(798), clk => clk, reset => reset); --
    end block;
    -- CP-element group 799:  join  transition  bypass 
    -- CP-element group 799: predecessors 
    -- CP-element group 799: 	792 
    -- CP-element group 799: 	795 
    -- CP-element group 799: 	798 
    -- CP-element group 799: successors 
    -- CP-element group 799: 	810 
    -- CP-element group 799:  members (1) 
      -- CP-element group 799: 	 branch_block_stmt_223/ifx_xelse1088_ifx_xend1126_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_799: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_799"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(792) & zeropad3D_CP_676_elements(795) & zeropad3D_CP_676_elements(798);
      gj_zeropad3D_cp_element_group_799 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(799), clk => clk, reset => reset); --
    end block;
    -- CP-element group 800:  transition  input  bypass 
    -- CP-element group 800: predecessors 
    -- CP-element group 800: 	387 
    -- CP-element group 800: successors 
    -- CP-element group 800: 	802 
    -- CP-element group 800:  members (2) 
      -- CP-element group 800: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Sample/$exit
      -- CP-element group 800: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Sample/ra
      -- 
    ra_8317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 800_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2607_inst_ack_0, ack => zeropad3D_CP_676_elements(800)); -- 
    -- CP-element group 801:  transition  input  bypass 
    -- CP-element group 801: predecessors 
    -- CP-element group 801: 	387 
    -- CP-element group 801: successors 
    -- CP-element group 801: 	802 
    -- CP-element group 801:  members (2) 
      -- CP-element group 801: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Update/$exit
      -- CP-element group 801: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/Update/ca
      -- 
    ca_8322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 801_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2607_inst_ack_1, ack => zeropad3D_CP_676_elements(801)); -- 
    -- CP-element group 802:  join  transition  output  bypass 
    -- CP-element group 802: predecessors 
    -- CP-element group 802: 	800 
    -- CP-element group 802: 	801 
    -- CP-element group 802: successors 
    -- CP-element group 802: 	809 
    -- CP-element group 802:  members (5) 
      -- CP-element group 802: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/$exit
      -- CP-element group 802: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/$exit
      -- CP-element group 802: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/$exit
      -- CP-element group 802: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_sources/type_cast_2607/SplitProtocol/$exit
      -- CP-element group 802: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2604/phi_stmt_2604_req
      -- 
    phi_stmt_2604_req_8323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2604_req_8323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(802), ack => phi_stmt_2604_req_0); -- 
    zeropad3D_cp_element_group_802: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_802"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(800) & zeropad3D_CP_676_elements(801);
      gj_zeropad3D_cp_element_group_802 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(802), clk => clk, reset => reset); --
    end block;
    -- CP-element group 803:  transition  input  bypass 
    -- CP-element group 803: predecessors 
    -- CP-element group 803: 	387 
    -- CP-element group 803: successors 
    -- CP-element group 803: 	805 
    -- CP-element group 803:  members (2) 
      -- CP-element group 803: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/SplitProtocol/Sample/$exit
      -- CP-element group 803: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/SplitProtocol/Sample/ra
      -- 
    ra_8340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 803_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_0, ack => zeropad3D_CP_676_elements(803)); -- 
    -- CP-element group 804:  transition  input  bypass 
    -- CP-element group 804: predecessors 
    -- CP-element group 804: 	387 
    -- CP-element group 804: successors 
    -- CP-element group 804: 	805 
    -- CP-element group 804:  members (2) 
      -- CP-element group 804: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/SplitProtocol/Update/$exit
      -- CP-element group 804: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/SplitProtocol/Update/ca
      -- 
    ca_8345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 804_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_1, ack => zeropad3D_CP_676_elements(804)); -- 
    -- CP-element group 805:  join  transition  output  bypass 
    -- CP-element group 805: predecessors 
    -- CP-element group 805: 	803 
    -- CP-element group 805: 	804 
    -- CP-element group 805: successors 
    -- CP-element group 805: 	809 
    -- CP-element group 805:  members (5) 
      -- CP-element group 805: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/$exit
      -- CP-element group 805: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/$exit
      -- CP-element group 805: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/$exit
      -- CP-element group 805: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_sources/type_cast_2614/SplitProtocol/$exit
      -- CP-element group 805: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2611/phi_stmt_2611_req
      -- 
    phi_stmt_2611_req_8346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2611_req_8346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(805), ack => phi_stmt_2611_req_0); -- 
    zeropad3D_cp_element_group_805: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_805"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(803) & zeropad3D_CP_676_elements(804);
      gj_zeropad3D_cp_element_group_805 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(805), clk => clk, reset => reset); --
    end block;
    -- CP-element group 806:  transition  input  bypass 
    -- CP-element group 806: predecessors 
    -- CP-element group 806: 	387 
    -- CP-element group 806: successors 
    -- CP-element group 806: 	808 
    -- CP-element group 806:  members (2) 
      -- CP-element group 806: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/SplitProtocol/Sample/$exit
      -- CP-element group 806: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/SplitProtocol/Sample/ra
      -- 
    ra_8363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 806_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2620_inst_ack_0, ack => zeropad3D_CP_676_elements(806)); -- 
    -- CP-element group 807:  transition  input  bypass 
    -- CP-element group 807: predecessors 
    -- CP-element group 807: 	387 
    -- CP-element group 807: successors 
    -- CP-element group 807: 	808 
    -- CP-element group 807:  members (2) 
      -- CP-element group 807: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/SplitProtocol/Update/$exit
      -- CP-element group 807: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/SplitProtocol/Update/ca
      -- 
    ca_8368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 807_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2620_inst_ack_1, ack => zeropad3D_CP_676_elements(807)); -- 
    -- CP-element group 808:  join  transition  output  bypass 
    -- CP-element group 808: predecessors 
    -- CP-element group 808: 	806 
    -- CP-element group 808: 	807 
    -- CP-element group 808: successors 
    -- CP-element group 808: 	809 
    -- CP-element group 808:  members (5) 
      -- CP-element group 808: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/$exit
      -- CP-element group 808: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/$exit
      -- CP-element group 808: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/$exit
      -- CP-element group 808: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_sources/type_cast_2620/SplitProtocol/$exit
      -- CP-element group 808: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/phi_stmt_2617/phi_stmt_2617_req
      -- 
    phi_stmt_2617_req_8369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2617_req_8369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(808), ack => phi_stmt_2617_req_0); -- 
    zeropad3D_cp_element_group_808: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_808"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(806) & zeropad3D_CP_676_elements(807);
      gj_zeropad3D_cp_element_group_808 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(808), clk => clk, reset => reset); --
    end block;
    -- CP-element group 809:  join  transition  bypass 
    -- CP-element group 809: predecessors 
    -- CP-element group 809: 	802 
    -- CP-element group 809: 	805 
    -- CP-element group 809: 	808 
    -- CP-element group 809: successors 
    -- CP-element group 809: 	810 
    -- CP-element group 809:  members (1) 
      -- CP-element group 809: 	 branch_block_stmt_223/ifx_xthen1083_ifx_xend1126_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_809: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_809"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(802) & zeropad3D_CP_676_elements(805) & zeropad3D_CP_676_elements(808);
      gj_zeropad3D_cp_element_group_809 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(809), clk => clk, reset => reset); --
    end block;
    -- CP-element group 810:  merge  fork  transition  place  bypass 
    -- CP-element group 810: predecessors 
    -- CP-element group 810: 	799 
    -- CP-element group 810: 	809 
    -- CP-element group 810: successors 
    -- CP-element group 810: 	811 
    -- CP-element group 810: 	812 
    -- CP-element group 810: 	813 
    -- CP-element group 810:  members (2) 
      -- CP-element group 810: 	 branch_block_stmt_223/merge_stmt_2603_PhiReqMerge
      -- CP-element group 810: 	 branch_block_stmt_223/merge_stmt_2603_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(810) <= OrReduce(zeropad3D_CP_676_elements(799) & zeropad3D_CP_676_elements(809));
    -- CP-element group 811:  transition  input  bypass 
    -- CP-element group 811: predecessors 
    -- CP-element group 811: 	810 
    -- CP-element group 811: successors 
    -- CP-element group 811: 	814 
    -- CP-element group 811:  members (1) 
      -- CP-element group 811: 	 branch_block_stmt_223/merge_stmt_2603_PhiAck/phi_stmt_2604_ack
      -- 
    phi_stmt_2604_ack_8374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 811_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2604_ack_0, ack => zeropad3D_CP_676_elements(811)); -- 
    -- CP-element group 812:  transition  input  bypass 
    -- CP-element group 812: predecessors 
    -- CP-element group 812: 	810 
    -- CP-element group 812: successors 
    -- CP-element group 812: 	814 
    -- CP-element group 812:  members (1) 
      -- CP-element group 812: 	 branch_block_stmt_223/merge_stmt_2603_PhiAck/phi_stmt_2611_ack
      -- 
    phi_stmt_2611_ack_8375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 812_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2611_ack_0, ack => zeropad3D_CP_676_elements(812)); -- 
    -- CP-element group 813:  transition  input  bypass 
    -- CP-element group 813: predecessors 
    -- CP-element group 813: 	810 
    -- CP-element group 813: successors 
    -- CP-element group 813: 	814 
    -- CP-element group 813:  members (1) 
      -- CP-element group 813: 	 branch_block_stmt_223/merge_stmt_2603_PhiAck/phi_stmt_2617_ack
      -- 
    phi_stmt_2617_ack_8376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 813_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2617_ack_0, ack => zeropad3D_CP_676_elements(813)); -- 
    -- CP-element group 814:  join  transition  bypass 
    -- CP-element group 814: predecessors 
    -- CP-element group 814: 	811 
    -- CP-element group 814: 	812 
    -- CP-element group 814: 	813 
    -- CP-element group 814: successors 
    -- CP-element group 814: 	5 
    -- CP-element group 814:  members (1) 
      -- CP-element group 814: 	 branch_block_stmt_223/merge_stmt_2603_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_814: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_814"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(811) & zeropad3D_CP_676_elements(812) & zeropad3D_CP_676_elements(813);
      gj_zeropad3D_cp_element_group_814 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(814), clk => clk, reset => reset); --
    end block;
    -- CP-element group 815:  transition  input  bypass 
    -- CP-element group 815: predecessors 
    -- CP-element group 815: 	6 
    -- CP-element group 815: successors 
    -- CP-element group 815: 	817 
    -- CP-element group 815:  members (2) 
      -- CP-element group 815: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/SplitProtocol/Sample/$exit
      -- CP-element group 815: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/SplitProtocol/Sample/ra
      -- 
    ra_8404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 815_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2667_inst_ack_0, ack => zeropad3D_CP_676_elements(815)); -- 
    -- CP-element group 816:  transition  input  bypass 
    -- CP-element group 816: predecessors 
    -- CP-element group 816: 	6 
    -- CP-element group 816: successors 
    -- CP-element group 816: 	817 
    -- CP-element group 816:  members (2) 
      -- CP-element group 816: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/SplitProtocol/Update/$exit
      -- CP-element group 816: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/SplitProtocol/Update/ca
      -- 
    ca_8409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 816_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2667_inst_ack_1, ack => zeropad3D_CP_676_elements(816)); -- 
    -- CP-element group 817:  join  transition  output  bypass 
    -- CP-element group 817: predecessors 
    -- CP-element group 817: 	815 
    -- CP-element group 817: 	816 
    -- CP-element group 817: successors 
    -- CP-element group 817: 	824 
    -- CP-element group 817:  members (5) 
      -- CP-element group 817: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/$exit
      -- CP-element group 817: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/$exit
      -- CP-element group 817: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/$exit
      -- CP-element group 817: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2667/SplitProtocol/$exit
      -- CP-element group 817: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_req
      -- 
    phi_stmt_2661_req_8410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2661_req_8410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(817), ack => phi_stmt_2661_req_1); -- 
    zeropad3D_cp_element_group_817: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_817"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(815) & zeropad3D_CP_676_elements(816);
      gj_zeropad3D_cp_element_group_817 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(817), clk => clk, reset => reset); --
    end block;
    -- CP-element group 818:  transition  input  bypass 
    -- CP-element group 818: predecessors 
    -- CP-element group 818: 	6 
    -- CP-element group 818: successors 
    -- CP-element group 818: 	820 
    -- CP-element group 818:  members (2) 
      -- CP-element group 818: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/SplitProtocol/Sample/$exit
      -- CP-element group 818: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/SplitProtocol/Sample/ra
      -- 
    ra_8427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 818_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2673_inst_ack_0, ack => zeropad3D_CP_676_elements(818)); -- 
    -- CP-element group 819:  transition  input  bypass 
    -- CP-element group 819: predecessors 
    -- CP-element group 819: 	6 
    -- CP-element group 819: successors 
    -- CP-element group 819: 	820 
    -- CP-element group 819:  members (2) 
      -- CP-element group 819: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/SplitProtocol/Update/$exit
      -- CP-element group 819: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/SplitProtocol/Update/ca
      -- 
    ca_8432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 819_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2673_inst_ack_1, ack => zeropad3D_CP_676_elements(819)); -- 
    -- CP-element group 820:  join  transition  output  bypass 
    -- CP-element group 820: predecessors 
    -- CP-element group 820: 	818 
    -- CP-element group 820: 	819 
    -- CP-element group 820: successors 
    -- CP-element group 820: 	824 
    -- CP-element group 820:  members (5) 
      -- CP-element group 820: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/$exit
      -- CP-element group 820: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/$exit
      -- CP-element group 820: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/$exit
      -- CP-element group 820: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2673/SplitProtocol/$exit
      -- CP-element group 820: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_req
      -- 
    phi_stmt_2668_req_8433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2668_req_8433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(820), ack => phi_stmt_2668_req_1); -- 
    zeropad3D_cp_element_group_820: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_820"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(818) & zeropad3D_CP_676_elements(819);
      gj_zeropad3D_cp_element_group_820 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(820), clk => clk, reset => reset); --
    end block;
    -- CP-element group 821:  transition  input  bypass 
    -- CP-element group 821: predecessors 
    -- CP-element group 821: 	6 
    -- CP-element group 821: successors 
    -- CP-element group 821: 	823 
    -- CP-element group 821:  members (2) 
      -- CP-element group 821: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/SplitProtocol/Sample/$exit
      -- CP-element group 821: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/SplitProtocol/Sample/ra
      -- 
    ra_8450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 821_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2679_inst_ack_0, ack => zeropad3D_CP_676_elements(821)); -- 
    -- CP-element group 822:  transition  input  bypass 
    -- CP-element group 822: predecessors 
    -- CP-element group 822: 	6 
    -- CP-element group 822: successors 
    -- CP-element group 822: 	823 
    -- CP-element group 822:  members (2) 
      -- CP-element group 822: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/SplitProtocol/Update/$exit
      -- CP-element group 822: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/SplitProtocol/Update/ca
      -- 
    ca_8455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 822_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2679_inst_ack_1, ack => zeropad3D_CP_676_elements(822)); -- 
    -- CP-element group 823:  join  transition  output  bypass 
    -- CP-element group 823: predecessors 
    -- CP-element group 823: 	821 
    -- CP-element group 823: 	822 
    -- CP-element group 823: successors 
    -- CP-element group 823: 	824 
    -- CP-element group 823:  members (5) 
      -- CP-element group 823: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/$exit
      -- CP-element group 823: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/$exit
      -- CP-element group 823: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/$exit
      -- CP-element group 823: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2679/SplitProtocol/$exit
      -- CP-element group 823: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_req
      -- 
    phi_stmt_2674_req_8456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2674_req_8456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(823), ack => phi_stmt_2674_req_1); -- 
    zeropad3D_cp_element_group_823: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_823"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(821) & zeropad3D_CP_676_elements(822);
      gj_zeropad3D_cp_element_group_823 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(823), clk => clk, reset => reset); --
    end block;
    -- CP-element group 824:  join  transition  bypass 
    -- CP-element group 824: predecessors 
    -- CP-element group 824: 	817 
    -- CP-element group 824: 	820 
    -- CP-element group 824: 	823 
    -- CP-element group 824: successors 
    -- CP-element group 824: 	833 
    -- CP-element group 824:  members (1) 
      -- CP-element group 824: 	 branch_block_stmt_223/ifx_xend1348_whilex_xbody1191_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_824: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_824"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(817) & zeropad3D_CP_676_elements(820) & zeropad3D_CP_676_elements(823);
      gj_zeropad3D_cp_element_group_824 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(824), clk => clk, reset => reset); --
    end block;
    -- CP-element group 825:  transition  output  delay-element  bypass 
    -- CP-element group 825: predecessors 
    -- CP-element group 825: 	400 
    -- CP-element group 825: successors 
    -- CP-element group 825: 	832 
    -- CP-element group 825:  members (4) 
      -- CP-element group 825: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2661/$exit
      -- CP-element group 825: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/$exit
      -- CP-element group 825: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_sources/type_cast_2665_konst_delay_trans
      -- CP-element group 825: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2661/phi_stmt_2661_req
      -- 
    phi_stmt_2661_req_8467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2661_req_8467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(825), ack => phi_stmt_2661_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(825) is a control-delay.
    cp_element_825_delay: control_delay_element  generic map(name => " 825_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(400), ack => zeropad3D_CP_676_elements(825), clk => clk, reset =>reset);
    -- CP-element group 826:  transition  input  bypass 
    -- CP-element group 826: predecessors 
    -- CP-element group 826: 	400 
    -- CP-element group 826: successors 
    -- CP-element group 826: 	828 
    -- CP-element group 826:  members (2) 
      -- CP-element group 826: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/SplitProtocol/Sample/$exit
      -- CP-element group 826: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/SplitProtocol/Sample/ra
      -- 
    ra_8484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 826_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2671_inst_ack_0, ack => zeropad3D_CP_676_elements(826)); -- 
    -- CP-element group 827:  transition  input  bypass 
    -- CP-element group 827: predecessors 
    -- CP-element group 827: 	400 
    -- CP-element group 827: successors 
    -- CP-element group 827: 	828 
    -- CP-element group 827:  members (2) 
      -- CP-element group 827: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/SplitProtocol/Update/$exit
      -- CP-element group 827: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/SplitProtocol/Update/ca
      -- 
    ca_8489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 827_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2671_inst_ack_1, ack => zeropad3D_CP_676_elements(827)); -- 
    -- CP-element group 828:  join  transition  output  bypass 
    -- CP-element group 828: predecessors 
    -- CP-element group 828: 	826 
    -- CP-element group 828: 	827 
    -- CP-element group 828: successors 
    -- CP-element group 828: 	832 
    -- CP-element group 828:  members (5) 
      -- CP-element group 828: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/$exit
      -- CP-element group 828: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/$exit
      -- CP-element group 828: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/$exit
      -- CP-element group 828: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_sources/type_cast_2671/SplitProtocol/$exit
      -- CP-element group 828: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2668/phi_stmt_2668_req
      -- 
    phi_stmt_2668_req_8490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2668_req_8490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(828), ack => phi_stmt_2668_req_0); -- 
    zeropad3D_cp_element_group_828: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_828"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(826) & zeropad3D_CP_676_elements(827);
      gj_zeropad3D_cp_element_group_828 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(828), clk => clk, reset => reset); --
    end block;
    -- CP-element group 829:  transition  input  bypass 
    -- CP-element group 829: predecessors 
    -- CP-element group 829: 	400 
    -- CP-element group 829: successors 
    -- CP-element group 829: 	831 
    -- CP-element group 829:  members (2) 
      -- CP-element group 829: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/SplitProtocol/Sample/$exit
      -- CP-element group 829: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/SplitProtocol/Sample/ra
      -- 
    ra_8507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 829_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2677_inst_ack_0, ack => zeropad3D_CP_676_elements(829)); -- 
    -- CP-element group 830:  transition  input  bypass 
    -- CP-element group 830: predecessors 
    -- CP-element group 830: 	400 
    -- CP-element group 830: successors 
    -- CP-element group 830: 	831 
    -- CP-element group 830:  members (2) 
      -- CP-element group 830: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/SplitProtocol/Update/$exit
      -- CP-element group 830: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/SplitProtocol/Update/ca
      -- 
    ca_8512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 830_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2677_inst_ack_1, ack => zeropad3D_CP_676_elements(830)); -- 
    -- CP-element group 831:  join  transition  output  bypass 
    -- CP-element group 831: predecessors 
    -- CP-element group 831: 	829 
    -- CP-element group 831: 	830 
    -- CP-element group 831: successors 
    -- CP-element group 831: 	832 
    -- CP-element group 831:  members (5) 
      -- CP-element group 831: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/$exit
      -- CP-element group 831: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/$exit
      -- CP-element group 831: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/$exit
      -- CP-element group 831: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_sources/type_cast_2677/SplitProtocol/$exit
      -- CP-element group 831: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/phi_stmt_2674/phi_stmt_2674_req
      -- 
    phi_stmt_2674_req_8513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2674_req_8513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(831), ack => phi_stmt_2674_req_0); -- 
    zeropad3D_cp_element_group_831: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_831"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(829) & zeropad3D_CP_676_elements(830);
      gj_zeropad3D_cp_element_group_831 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(831), clk => clk, reset => reset); --
    end block;
    -- CP-element group 832:  join  transition  bypass 
    -- CP-element group 832: predecessors 
    -- CP-element group 832: 	825 
    -- CP-element group 832: 	828 
    -- CP-element group 832: 	831 
    -- CP-element group 832: successors 
    -- CP-element group 832: 	833 
    -- CP-element group 832:  members (1) 
      -- CP-element group 832: 	 branch_block_stmt_223/whilex_xend1127_whilex_xbody1191_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_832: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_832"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(825) & zeropad3D_CP_676_elements(828) & zeropad3D_CP_676_elements(831);
      gj_zeropad3D_cp_element_group_832 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(832), clk => clk, reset => reset); --
    end block;
    -- CP-element group 833:  merge  fork  transition  place  bypass 
    -- CP-element group 833: predecessors 
    -- CP-element group 833: 	824 
    -- CP-element group 833: 	832 
    -- CP-element group 833: successors 
    -- CP-element group 833: 	834 
    -- CP-element group 833: 	835 
    -- CP-element group 833: 	836 
    -- CP-element group 833:  members (2) 
      -- CP-element group 833: 	 branch_block_stmt_223/merge_stmt_2660_PhiReqMerge
      -- CP-element group 833: 	 branch_block_stmt_223/merge_stmt_2660_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(833) <= OrReduce(zeropad3D_CP_676_elements(824) & zeropad3D_CP_676_elements(832));
    -- CP-element group 834:  transition  input  bypass 
    -- CP-element group 834: predecessors 
    -- CP-element group 834: 	833 
    -- CP-element group 834: successors 
    -- CP-element group 834: 	837 
    -- CP-element group 834:  members (1) 
      -- CP-element group 834: 	 branch_block_stmt_223/merge_stmt_2660_PhiAck/phi_stmt_2661_ack
      -- 
    phi_stmt_2661_ack_8518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 834_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2661_ack_0, ack => zeropad3D_CP_676_elements(834)); -- 
    -- CP-element group 835:  transition  input  bypass 
    -- CP-element group 835: predecessors 
    -- CP-element group 835: 	833 
    -- CP-element group 835: successors 
    -- CP-element group 835: 	837 
    -- CP-element group 835:  members (1) 
      -- CP-element group 835: 	 branch_block_stmt_223/merge_stmt_2660_PhiAck/phi_stmt_2668_ack
      -- 
    phi_stmt_2668_ack_8519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 835_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2668_ack_0, ack => zeropad3D_CP_676_elements(835)); -- 
    -- CP-element group 836:  transition  input  bypass 
    -- CP-element group 836: predecessors 
    -- CP-element group 836: 	833 
    -- CP-element group 836: successors 
    -- CP-element group 836: 	837 
    -- CP-element group 836:  members (1) 
      -- CP-element group 836: 	 branch_block_stmt_223/merge_stmt_2660_PhiAck/phi_stmt_2674_ack
      -- 
    phi_stmt_2674_ack_8520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 836_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2674_ack_0, ack => zeropad3D_CP_676_elements(836)); -- 
    -- CP-element group 837:  join  fork  transition  place  output  bypass 
    -- CP-element group 837: predecessors 
    -- CP-element group 837: 	834 
    -- CP-element group 837: 	835 
    -- CP-element group 837: 	836 
    -- CP-element group 837: successors 
    -- CP-element group 837: 	401 
    -- CP-element group 837: 	402 
    -- CP-element group 837:  members (10) 
      -- CP-element group 837: 	 branch_block_stmt_223/merge_stmt_2660__exit__
      -- CP-element group 837: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710__entry__
      -- CP-element group 837: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/$entry
      -- CP-element group 837: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_sample_start_
      -- CP-element group 837: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_update_start_
      -- CP-element group 837: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_Sample/$entry
      -- CP-element group 837: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_Sample/rr
      -- CP-element group 837: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_Update/$entry
      -- CP-element group 837: 	 branch_block_stmt_223/assign_stmt_2685_to_assign_stmt_2710/type_cast_2684_Update/cr
      -- CP-element group 837: 	 branch_block_stmt_223/merge_stmt_2660_PhiAck/$exit
      -- 
    rr_4839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(837), ack => type_cast_2684_inst_req_0); -- 
    cr_4844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(837), ack => type_cast_2684_inst_req_1); -- 
    zeropad3D_cp_element_group_837: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_837"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(834) & zeropad3D_CP_676_elements(835) & zeropad3D_CP_676_elements(836);
      gj_zeropad3D_cp_element_group_837 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(837), clk => clk, reset => reset); --
    end block;
    -- CP-element group 838:  merge  fork  transition  place  output  bypass 
    -- CP-element group 838: predecessors 
    -- CP-element group 838: 	404 
    -- CP-element group 838: 	408 
    -- CP-element group 838: successors 
    -- CP-element group 838: 	409 
    -- CP-element group 838: 	410 
    -- CP-element group 838: 	411 
    -- CP-element group 838: 	412 
    -- CP-element group 838: 	415 
    -- CP-element group 838: 	417 
    -- CP-element group 838: 	419 
    -- CP-element group 838: 	421 
    -- CP-element group 838:  members (33) 
      -- CP-element group 838: 	 branch_block_stmt_223/merge_stmt_2754__exit__
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810__entry__
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Update/word_access_complete/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_complete/req
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_update_start_
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_Update/cr
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Update/word_access_complete/word_0/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_update_start_
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_final_index_sum_regn_update_start
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Update/word_access_complete/word_0/cr
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_update_start_
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_final_index_sum_regn_Update/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/array_obj_ref_2803_final_index_sum_regn_Update/req
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/ptr_deref_2807_Update/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_Update/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/addr_of_2804_complete/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_Sample/rr
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_Update/cr
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2797_Update/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_sample_start_
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_update_start_
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_Sample/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_Sample/rr
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_Update/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2758_Update/cr
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_sample_start_
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_update_start_
      -- CP-element group 838: 	 branch_block_stmt_223/assign_stmt_2759_to_assign_stmt_2810/type_cast_2763_Sample/$entry
      -- CP-element group 838: 	 branch_block_stmt_223/merge_stmt_2754_PhiReqMerge
      -- CP-element group 838: 	 branch_block_stmt_223/merge_stmt_2754_PhiAck/dummy
      -- CP-element group 838: 	 branch_block_stmt_223/merge_stmt_2754_PhiAck/$exit
      -- CP-element group 838: 	 branch_block_stmt_223/merge_stmt_2754_PhiAck/$entry
      -- 
    req_4990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(838), ack => addr_of_2804_final_reg_req_1); -- 
    cr_4930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(838), ack => type_cast_2763_inst_req_1); -- 
    cr_5040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(838), ack => ptr_deref_2807_store_0_req_1); -- 
    req_4975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(838), ack => array_obj_ref_2803_index_offset_req_1); -- 
    rr_4925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(838), ack => type_cast_2763_inst_req_0); -- 
    cr_4944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(838), ack => type_cast_2797_inst_req_1); -- 
    rr_4911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(838), ack => type_cast_2758_inst_req_0); -- 
    cr_4916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(838), ack => type_cast_2758_inst_req_1); -- 
    zeropad3D_CP_676_elements(838) <= OrReduce(zeropad3D_CP_676_elements(404) & zeropad3D_CP_676_elements(408));
    -- CP-element group 839:  merge  fork  transition  place  output  bypass 
    -- CP-element group 839: predecessors 
    -- CP-element group 839: 	422 
    -- CP-element group 839: 	442 
    -- CP-element group 839: successors 
    -- CP-element group 839: 	443 
    -- CP-element group 839: 	444 
    -- CP-element group 839:  members (13) 
      -- CP-element group 839: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937__entry__
      -- CP-element group 839: 	 branch_block_stmt_223/merge_stmt_2919__exit__
      -- CP-element group 839: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/$entry
      -- CP-element group 839: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_sample_start_
      -- CP-element group 839: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_update_start_
      -- CP-element group 839: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_Sample/$entry
      -- CP-element group 839: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_Sample/rr
      -- CP-element group 839: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_Update/$entry
      -- CP-element group 839: 	 branch_block_stmt_223/assign_stmt_2924_to_assign_stmt_2937/type_cast_2923_Update/cr
      -- CP-element group 839: 	 branch_block_stmt_223/merge_stmt_2919_PhiAck/dummy
      -- CP-element group 839: 	 branch_block_stmt_223/merge_stmt_2919_PhiAck/$exit
      -- CP-element group 839: 	 branch_block_stmt_223/merge_stmt_2919_PhiAck/$entry
      -- CP-element group 839: 	 branch_block_stmt_223/merge_stmt_2919_PhiReqMerge
      -- 
    rr_5289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(839), ack => type_cast_2923_inst_req_0); -- 
    cr_5294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(839), ack => type_cast_2923_inst_req_1); -- 
    zeropad3D_CP_676_elements(839) <= OrReduce(zeropad3D_CP_676_elements(422) & zeropad3D_CP_676_elements(442));
    -- CP-element group 840:  transition  output  delay-element  bypass 
    -- CP-element group 840: predecessors 
    -- CP-element group 840: 	454 
    -- CP-element group 840: successors 
    -- CP-element group 840: 	847 
    -- CP-element group 840:  members (4) 
      -- CP-element group 840: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_req
      -- CP-element group 840: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3007_konst_delay_trans
      -- CP-element group 840: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/$exit
      -- CP-element group 840: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3001/$exit
      -- 
    phi_stmt_3001_req_8601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3001_req_8601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(840), ack => phi_stmt_3001_req_1); -- 
    -- Element group zeropad3D_CP_676_elements(840) is a control-delay.
    cp_element_840_delay: control_delay_element  generic map(name => " 840_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(454), ack => zeropad3D_CP_676_elements(840), clk => clk, reset =>reset);
    -- CP-element group 841:  transition  input  bypass 
    -- CP-element group 841: predecessors 
    -- CP-element group 841: 	454 
    -- CP-element group 841: successors 
    -- CP-element group 841: 	843 
    -- CP-element group 841:  members (2) 
      -- CP-element group 841: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/SplitProtocol/Sample/ra
      -- CP-element group 841: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/SplitProtocol/Sample/$exit
      -- 
    ra_8618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 841_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3013_inst_ack_0, ack => zeropad3D_CP_676_elements(841)); -- 
    -- CP-element group 842:  transition  input  bypass 
    -- CP-element group 842: predecessors 
    -- CP-element group 842: 	454 
    -- CP-element group 842: successors 
    -- CP-element group 842: 	843 
    -- CP-element group 842:  members (2) 
      -- CP-element group 842: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/SplitProtocol/Update/ca
      -- CP-element group 842: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/SplitProtocol/Update/$exit
      -- 
    ca_8623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 842_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3013_inst_ack_1, ack => zeropad3D_CP_676_elements(842)); -- 
    -- CP-element group 843:  join  transition  output  bypass 
    -- CP-element group 843: predecessors 
    -- CP-element group 843: 	841 
    -- CP-element group 843: 	842 
    -- CP-element group 843: successors 
    -- CP-element group 843: 	847 
    -- CP-element group 843:  members (5) 
      -- CP-element group 843: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/$exit
      -- CP-element group 843: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/$exit
      -- CP-element group 843: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/$exit
      -- CP-element group 843: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3013/SplitProtocol/$exit
      -- CP-element group 843: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_req
      -- 
    phi_stmt_3008_req_8624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3008_req_8624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(843), ack => phi_stmt_3008_req_1); -- 
    zeropad3D_cp_element_group_843: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_843"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(841) & zeropad3D_CP_676_elements(842);
      gj_zeropad3D_cp_element_group_843 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(843), clk => clk, reset => reset); --
    end block;
    -- CP-element group 844:  transition  input  bypass 
    -- CP-element group 844: predecessors 
    -- CP-element group 844: 	454 
    -- CP-element group 844: successors 
    -- CP-element group 844: 	846 
    -- CP-element group 844:  members (2) 
      -- CP-element group 844: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/SplitProtocol/Sample/$exit
      -- CP-element group 844: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/SplitProtocol/Sample/ra
      -- 
    ra_8641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 844_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3019_inst_ack_0, ack => zeropad3D_CP_676_elements(844)); -- 
    -- CP-element group 845:  transition  input  bypass 
    -- CP-element group 845: predecessors 
    -- CP-element group 845: 	454 
    -- CP-element group 845: successors 
    -- CP-element group 845: 	846 
    -- CP-element group 845:  members (2) 
      -- CP-element group 845: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/SplitProtocol/Update/ca
      -- CP-element group 845: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/SplitProtocol/Update/$exit
      -- 
    ca_8646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 845_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3019_inst_ack_1, ack => zeropad3D_CP_676_elements(845)); -- 
    -- CP-element group 846:  join  transition  output  bypass 
    -- CP-element group 846: predecessors 
    -- CP-element group 846: 	844 
    -- CP-element group 846: 	845 
    -- CP-element group 846: successors 
    -- CP-element group 846: 	847 
    -- CP-element group 846:  members (5) 
      -- CP-element group 846: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/SplitProtocol/$exit
      -- CP-element group 846: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3019/$exit
      -- CP-element group 846: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/$exit
      -- CP-element group 846: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/$exit
      -- CP-element group 846: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_req
      -- 
    phi_stmt_3014_req_8647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3014_req_8647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(846), ack => phi_stmt_3014_req_1); -- 
    zeropad3D_cp_element_group_846: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_846"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(844) & zeropad3D_CP_676_elements(845);
      gj_zeropad3D_cp_element_group_846 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(846), clk => clk, reset => reset); --
    end block;
    -- CP-element group 847:  join  transition  bypass 
    -- CP-element group 847: predecessors 
    -- CP-element group 847: 	840 
    -- CP-element group 847: 	843 
    -- CP-element group 847: 	846 
    -- CP-element group 847: successors 
    -- CP-element group 847: 	858 
    -- CP-element group 847:  members (1) 
      -- CP-element group 847: 	 branch_block_stmt_223/ifx_xelse1311_ifx_xend1348_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_847: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_847"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(840) & zeropad3D_CP_676_elements(843) & zeropad3D_CP_676_elements(846);
      gj_zeropad3D_cp_element_group_847 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(847), clk => clk, reset => reset); --
    end block;
    -- CP-element group 848:  transition  input  bypass 
    -- CP-element group 848: predecessors 
    -- CP-element group 848: 	445 
    -- CP-element group 848: successors 
    -- CP-element group 848: 	850 
    -- CP-element group 848:  members (2) 
      -- CP-element group 848: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/SplitProtocol/Sample/ra
      -- CP-element group 848: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/SplitProtocol/Sample/$exit
      -- 
    ra_8667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 848_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3004_inst_ack_0, ack => zeropad3D_CP_676_elements(848)); -- 
    -- CP-element group 849:  transition  input  bypass 
    -- CP-element group 849: predecessors 
    -- CP-element group 849: 	445 
    -- CP-element group 849: successors 
    -- CP-element group 849: 	850 
    -- CP-element group 849:  members (2) 
      -- CP-element group 849: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/SplitProtocol/Update/ca
      -- CP-element group 849: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/SplitProtocol/Update/$exit
      -- 
    ca_8672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 849_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3004_inst_ack_1, ack => zeropad3D_CP_676_elements(849)); -- 
    -- CP-element group 850:  join  transition  output  bypass 
    -- CP-element group 850: predecessors 
    -- CP-element group 850: 	848 
    -- CP-element group 850: 	849 
    -- CP-element group 850: successors 
    -- CP-element group 850: 	857 
    -- CP-element group 850:  members (5) 
      -- CP-element group 850: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_req
      -- CP-element group 850: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/SplitProtocol/$exit
      -- CP-element group 850: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/type_cast_3004/$exit
      -- CP-element group 850: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/phi_stmt_3001_sources/$exit
      -- CP-element group 850: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3001/$exit
      -- 
    phi_stmt_3001_req_8673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3001_req_8673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(850), ack => phi_stmt_3001_req_0); -- 
    zeropad3D_cp_element_group_850: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_850"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(848) & zeropad3D_CP_676_elements(849);
      gj_zeropad3D_cp_element_group_850 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(850), clk => clk, reset => reset); --
    end block;
    -- CP-element group 851:  transition  input  bypass 
    -- CP-element group 851: predecessors 
    -- CP-element group 851: 	445 
    -- CP-element group 851: successors 
    -- CP-element group 851: 	853 
    -- CP-element group 851:  members (2) 
      -- CP-element group 851: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/SplitProtocol/Sample/$exit
      -- CP-element group 851: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/SplitProtocol/Sample/ra
      -- 
    ra_8690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 851_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3011_inst_ack_0, ack => zeropad3D_CP_676_elements(851)); -- 
    -- CP-element group 852:  transition  input  bypass 
    -- CP-element group 852: predecessors 
    -- CP-element group 852: 	445 
    -- CP-element group 852: successors 
    -- CP-element group 852: 	853 
    -- CP-element group 852:  members (2) 
      -- CP-element group 852: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/SplitProtocol/Update/ca
      -- CP-element group 852: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/SplitProtocol/Update/$exit
      -- 
    ca_8695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 852_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3011_inst_ack_1, ack => zeropad3D_CP_676_elements(852)); -- 
    -- CP-element group 853:  join  transition  output  bypass 
    -- CP-element group 853: predecessors 
    -- CP-element group 853: 	851 
    -- CP-element group 853: 	852 
    -- CP-element group 853: successors 
    -- CP-element group 853: 	857 
    -- CP-element group 853:  members (5) 
      -- CP-element group 853: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/$exit
      -- CP-element group 853: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/$exit
      -- CP-element group 853: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/$exit
      -- CP-element group 853: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_sources/type_cast_3011/SplitProtocol/$exit
      -- CP-element group 853: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3008/phi_stmt_3008_req
      -- 
    phi_stmt_3008_req_8696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3008_req_8696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(853), ack => phi_stmt_3008_req_0); -- 
    zeropad3D_cp_element_group_853: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_853"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(851) & zeropad3D_CP_676_elements(852);
      gj_zeropad3D_cp_element_group_853 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(853), clk => clk, reset => reset); --
    end block;
    -- CP-element group 854:  transition  input  bypass 
    -- CP-element group 854: predecessors 
    -- CP-element group 854: 	445 
    -- CP-element group 854: successors 
    -- CP-element group 854: 	856 
    -- CP-element group 854:  members (2) 
      -- CP-element group 854: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/SplitProtocol/Sample/ra
      -- CP-element group 854: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/SplitProtocol/Sample/$exit
      -- 
    ra_8713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 854_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3017_inst_ack_0, ack => zeropad3D_CP_676_elements(854)); -- 
    -- CP-element group 855:  transition  input  bypass 
    -- CP-element group 855: predecessors 
    -- CP-element group 855: 	445 
    -- CP-element group 855: successors 
    -- CP-element group 855: 	856 
    -- CP-element group 855:  members (2) 
      -- CP-element group 855: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/SplitProtocol/Update/ca
      -- CP-element group 855: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/SplitProtocol/Update/$exit
      -- 
    ca_8718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 855_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3017_inst_ack_1, ack => zeropad3D_CP_676_elements(855)); -- 
    -- CP-element group 856:  join  transition  output  bypass 
    -- CP-element group 856: predecessors 
    -- CP-element group 856: 	854 
    -- CP-element group 856: 	855 
    -- CP-element group 856: successors 
    -- CP-element group 856: 	857 
    -- CP-element group 856:  members (5) 
      -- CP-element group 856: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/$exit
      -- CP-element group 856: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_req
      -- CP-element group 856: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/SplitProtocol/$exit
      -- CP-element group 856: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/type_cast_3017/$exit
      -- CP-element group 856: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/phi_stmt_3014/phi_stmt_3014_sources/$exit
      -- 
    phi_stmt_3014_req_8719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3014_req_8719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(856), ack => phi_stmt_3014_req_0); -- 
    zeropad3D_cp_element_group_856: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_856"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(854) & zeropad3D_CP_676_elements(855);
      gj_zeropad3D_cp_element_group_856 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(856), clk => clk, reset => reset); --
    end block;
    -- CP-element group 857:  join  transition  bypass 
    -- CP-element group 857: predecessors 
    -- CP-element group 857: 	850 
    -- CP-element group 857: 	853 
    -- CP-element group 857: 	856 
    -- CP-element group 857: successors 
    -- CP-element group 857: 	858 
    -- CP-element group 857:  members (1) 
      -- CP-element group 857: 	 branch_block_stmt_223/ifx_xthen1306_ifx_xend1348_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_857: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_857"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(850) & zeropad3D_CP_676_elements(853) & zeropad3D_CP_676_elements(856);
      gj_zeropad3D_cp_element_group_857 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(857), clk => clk, reset => reset); --
    end block;
    -- CP-element group 858:  merge  fork  transition  place  bypass 
    -- CP-element group 858: predecessors 
    -- CP-element group 858: 	847 
    -- CP-element group 858: 	857 
    -- CP-element group 858: successors 
    -- CP-element group 858: 	859 
    -- CP-element group 858: 	860 
    -- CP-element group 858: 	861 
    -- CP-element group 858:  members (2) 
      -- CP-element group 858: 	 branch_block_stmt_223/merge_stmt_3000_PhiAck/$entry
      -- CP-element group 858: 	 branch_block_stmt_223/merge_stmt_3000_PhiReqMerge
      -- 
    zeropad3D_CP_676_elements(858) <= OrReduce(zeropad3D_CP_676_elements(847) & zeropad3D_CP_676_elements(857));
    -- CP-element group 859:  transition  input  bypass 
    -- CP-element group 859: predecessors 
    -- CP-element group 859: 	858 
    -- CP-element group 859: successors 
    -- CP-element group 859: 	862 
    -- CP-element group 859:  members (1) 
      -- CP-element group 859: 	 branch_block_stmt_223/merge_stmt_3000_PhiAck/phi_stmt_3001_ack
      -- 
    phi_stmt_3001_ack_8724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 859_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3001_ack_0, ack => zeropad3D_CP_676_elements(859)); -- 
    -- CP-element group 860:  transition  input  bypass 
    -- CP-element group 860: predecessors 
    -- CP-element group 860: 	858 
    -- CP-element group 860: successors 
    -- CP-element group 860: 	862 
    -- CP-element group 860:  members (1) 
      -- CP-element group 860: 	 branch_block_stmt_223/merge_stmt_3000_PhiAck/phi_stmt_3008_ack
      -- 
    phi_stmt_3008_ack_8725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 860_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3008_ack_0, ack => zeropad3D_CP_676_elements(860)); -- 
    -- CP-element group 861:  transition  input  bypass 
    -- CP-element group 861: predecessors 
    -- CP-element group 861: 	858 
    -- CP-element group 861: successors 
    -- CP-element group 861: 	862 
    -- CP-element group 861:  members (1) 
      -- CP-element group 861: 	 branch_block_stmt_223/merge_stmt_3000_PhiAck/phi_stmt_3014_ack
      -- 
    phi_stmt_3014_ack_8726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 861_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3014_ack_0, ack => zeropad3D_CP_676_elements(861)); -- 
    -- CP-element group 862:  join  transition  bypass 
    -- CP-element group 862: predecessors 
    -- CP-element group 862: 	859 
    -- CP-element group 862: 	860 
    -- CP-element group 862: 	861 
    -- CP-element group 862: successors 
    -- CP-element group 862: 	6 
    -- CP-element group 862:  members (1) 
      -- CP-element group 862: 	 branch_block_stmt_223/merge_stmt_3000_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_862: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_862"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(859) & zeropad3D_CP_676_elements(860) & zeropad3D_CP_676_elements(861);
      gj_zeropad3D_cp_element_group_862 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(862), clk => clk, reset => reset); --
    end block;
    -- CP-element group 863:  transition  input  bypass 
    -- CP-element group 863: predecessors 
    -- CP-element group 863: 	7 
    -- CP-element group 863: successors 
    -- CP-element group 863: 	865 
    -- CP-element group 863:  members (2) 
      -- CP-element group 863: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/SplitProtocol/Sample/ra
      -- CP-element group 863: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/SplitProtocol/Sample/$exit
      -- 
    ra_8754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 863_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3080_inst_ack_0, ack => zeropad3D_CP_676_elements(863)); -- 
    -- CP-element group 864:  transition  input  bypass 
    -- CP-element group 864: predecessors 
    -- CP-element group 864: 	7 
    -- CP-element group 864: successors 
    -- CP-element group 864: 	865 
    -- CP-element group 864:  members (2) 
      -- CP-element group 864: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/SplitProtocol/Update/$exit
      -- CP-element group 864: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/SplitProtocol/Update/ca
      -- 
    ca_8759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 864_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3080_inst_ack_1, ack => zeropad3D_CP_676_elements(864)); -- 
    -- CP-element group 865:  join  transition  output  bypass 
    -- CP-element group 865: predecessors 
    -- CP-element group 865: 	863 
    -- CP-element group 865: 	864 
    -- CP-element group 865: successors 
    -- CP-element group 865: 	872 
    -- CP-element group 865:  members (5) 
      -- CP-element group 865: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/$exit
      -- CP-element group 865: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/$exit
      -- CP-element group 865: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/SplitProtocol/$exit
      -- CP-element group 865: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_req
      -- CP-element group 865: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3080/$exit
      -- 
    phi_stmt_3077_req_8760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3077_req_8760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(865), ack => phi_stmt_3077_req_0); -- 
    zeropad3D_cp_element_group_865: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_865"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(863) & zeropad3D_CP_676_elements(864);
      gj_zeropad3D_cp_element_group_865 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(865), clk => clk, reset => reset); --
    end block;
    -- CP-element group 866:  transition  input  bypass 
    -- CP-element group 866: predecessors 
    -- CP-element group 866: 	7 
    -- CP-element group 866: successors 
    -- CP-element group 866: 	868 
    -- CP-element group 866:  members (2) 
      -- CP-element group 866: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/SplitProtocol/Sample/ra
      -- CP-element group 866: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/SplitProtocol/Sample/$exit
      -- 
    ra_8777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 866_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3070_inst_ack_0, ack => zeropad3D_CP_676_elements(866)); -- 
    -- CP-element group 867:  transition  input  bypass 
    -- CP-element group 867: predecessors 
    -- CP-element group 867: 	7 
    -- CP-element group 867: successors 
    -- CP-element group 867: 	868 
    -- CP-element group 867:  members (2) 
      -- CP-element group 867: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/SplitProtocol/Update/ca
      -- CP-element group 867: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/SplitProtocol/Update/$exit
      -- 
    ca_8782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 867_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3070_inst_ack_1, ack => zeropad3D_CP_676_elements(867)); -- 
    -- CP-element group 868:  join  transition  output  bypass 
    -- CP-element group 868: predecessors 
    -- CP-element group 868: 	866 
    -- CP-element group 868: 	867 
    -- CP-element group 868: successors 
    -- CP-element group 868: 	872 
    -- CP-element group 868:  members (5) 
      -- CP-element group 868: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/$exit
      -- CP-element group 868: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/$exit
      -- CP-element group 868: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/$exit
      -- CP-element group 868: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_req
      -- CP-element group 868: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3070/SplitProtocol/$exit
      -- 
    phi_stmt_3064_req_8783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3064_req_8783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(868), ack => phi_stmt_3064_req_1); -- 
    zeropad3D_cp_element_group_868: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_868"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(866) & zeropad3D_CP_676_elements(867);
      gj_zeropad3D_cp_element_group_868 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(868), clk => clk, reset => reset); --
    end block;
    -- CP-element group 869:  transition  input  bypass 
    -- CP-element group 869: predecessors 
    -- CP-element group 869: 	7 
    -- CP-element group 869: successors 
    -- CP-element group 869: 	871 
    -- CP-element group 869:  members (2) 
      -- CP-element group 869: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/SplitProtocol/Sample/ra
      -- CP-element group 869: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/SplitProtocol/Sample/$exit
      -- 
    ra_8800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 869_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3074_inst_ack_0, ack => zeropad3D_CP_676_elements(869)); -- 
    -- CP-element group 870:  transition  input  bypass 
    -- CP-element group 870: predecessors 
    -- CP-element group 870: 	7 
    -- CP-element group 870: successors 
    -- CP-element group 870: 	871 
    -- CP-element group 870:  members (2) 
      -- CP-element group 870: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/SplitProtocol/Update/ca
      -- CP-element group 870: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/SplitProtocol/Update/$exit
      -- 
    ca_8805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 870_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3074_inst_ack_1, ack => zeropad3D_CP_676_elements(870)); -- 
    -- CP-element group 871:  join  transition  output  bypass 
    -- CP-element group 871: predecessors 
    -- CP-element group 871: 	869 
    -- CP-element group 871: 	870 
    -- CP-element group 871: successors 
    -- CP-element group 871: 	872 
    -- CP-element group 871:  members (5) 
      -- CP-element group 871: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/SplitProtocol/$exit
      -- CP-element group 871: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_req
      -- CP-element group 871: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3074/$exit
      -- CP-element group 871: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/$exit
      -- CP-element group 871: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/phi_stmt_3071/$exit
      -- 
    phi_stmt_3071_req_8806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3071_req_8806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(871), ack => phi_stmt_3071_req_0); -- 
    zeropad3D_cp_element_group_871: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_871"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(869) & zeropad3D_CP_676_elements(870);
      gj_zeropad3D_cp_element_group_871 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(871), clk => clk, reset => reset); --
    end block;
    -- CP-element group 872:  join  transition  bypass 
    -- CP-element group 872: predecessors 
    -- CP-element group 872: 	865 
    -- CP-element group 872: 	868 
    -- CP-element group 872: 	871 
    -- CP-element group 872: successors 
    -- CP-element group 872: 	879 
    -- CP-element group 872:  members (1) 
      -- CP-element group 872: 	 branch_block_stmt_223/ifx_xend1565_whilex_xbody1410_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_872: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_872"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(865) & zeropad3D_CP_676_elements(868) & zeropad3D_CP_676_elements(871);
      gj_zeropad3D_cp_element_group_872 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(872), clk => clk, reset => reset); --
    end block;
    -- CP-element group 873:  transition  output  delay-element  bypass 
    -- CP-element group 873: predecessors 
    -- CP-element group 873: 	458 
    -- CP-element group 873: successors 
    -- CP-element group 873: 	878 
    -- CP-element group 873:  members (4) 
      -- CP-element group 873: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3077/$exit
      -- CP-element group 873: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/$exit
      -- CP-element group 873: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_sources/type_cast_3083_konst_delay_trans
      -- CP-element group 873: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3077/phi_stmt_3077_req
      -- 
    phi_stmt_3077_req_8817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3077_req_8817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(873), ack => phi_stmt_3077_req_1); -- 
    -- Element group zeropad3D_CP_676_elements(873) is a control-delay.
    cp_element_873_delay: control_delay_element  generic map(name => " 873_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(458), ack => zeropad3D_CP_676_elements(873), clk => clk, reset =>reset);
    -- CP-element group 874:  transition  output  delay-element  bypass 
    -- CP-element group 874: predecessors 
    -- CP-element group 874: 	458 
    -- CP-element group 874: successors 
    -- CP-element group 874: 	878 
    -- CP-element group 874:  members (4) 
      -- CP-element group 874: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3064/$exit
      -- CP-element group 874: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/$exit
      -- CP-element group 874: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_sources/type_cast_3068_konst_delay_trans
      -- CP-element group 874: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3064/phi_stmt_3064_req
      -- 
    phi_stmt_3064_req_8825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3064_req_8825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(874), ack => phi_stmt_3064_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(874) is a control-delay.
    cp_element_874_delay: control_delay_element  generic map(name => " 874_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(458), ack => zeropad3D_CP_676_elements(874), clk => clk, reset =>reset);
    -- CP-element group 875:  transition  input  bypass 
    -- CP-element group 875: predecessors 
    -- CP-element group 875: 	458 
    -- CP-element group 875: successors 
    -- CP-element group 875: 	877 
    -- CP-element group 875:  members (2) 
      -- CP-element group 875: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/SplitProtocol/Sample/$exit
      -- CP-element group 875: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/SplitProtocol/Sample/ra
      -- 
    ra_8842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 875_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3076_inst_ack_0, ack => zeropad3D_CP_676_elements(875)); -- 
    -- CP-element group 876:  transition  input  bypass 
    -- CP-element group 876: predecessors 
    -- CP-element group 876: 	458 
    -- CP-element group 876: successors 
    -- CP-element group 876: 	877 
    -- CP-element group 876:  members (2) 
      -- CP-element group 876: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/SplitProtocol/Update/$exit
      -- CP-element group 876: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/SplitProtocol/Update/ca
      -- 
    ca_8847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 876_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3076_inst_ack_1, ack => zeropad3D_CP_676_elements(876)); -- 
    -- CP-element group 877:  join  transition  output  bypass 
    -- CP-element group 877: predecessors 
    -- CP-element group 877: 	875 
    -- CP-element group 877: 	876 
    -- CP-element group 877: successors 
    -- CP-element group 877: 	878 
    -- CP-element group 877:  members (5) 
      -- CP-element group 877: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/$exit
      -- CP-element group 877: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/$exit
      -- CP-element group 877: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/$exit
      -- CP-element group 877: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_sources/type_cast_3076/SplitProtocol/$exit
      -- CP-element group 877: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/phi_stmt_3071/phi_stmt_3071_req
      -- 
    phi_stmt_3071_req_8848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3071_req_8848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(877), ack => phi_stmt_3071_req_1); -- 
    zeropad3D_cp_element_group_877: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_877"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(875) & zeropad3D_CP_676_elements(876);
      gj_zeropad3D_cp_element_group_877 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(877), clk => clk, reset => reset); --
    end block;
    -- CP-element group 878:  join  transition  bypass 
    -- CP-element group 878: predecessors 
    -- CP-element group 878: 	873 
    -- CP-element group 878: 	874 
    -- CP-element group 878: 	877 
    -- CP-element group 878: successors 
    -- CP-element group 878: 	879 
    -- CP-element group 878:  members (1) 
      -- CP-element group 878: 	 branch_block_stmt_223/whilex_xend1349_whilex_xbody1410_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_878: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_878"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(873) & zeropad3D_CP_676_elements(874) & zeropad3D_CP_676_elements(877);
      gj_zeropad3D_cp_element_group_878 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(878), clk => clk, reset => reset); --
    end block;
    -- CP-element group 879:  merge  fork  transition  place  bypass 
    -- CP-element group 879: predecessors 
    -- CP-element group 879: 	872 
    -- CP-element group 879: 	878 
    -- CP-element group 879: successors 
    -- CP-element group 879: 	880 
    -- CP-element group 879: 	881 
    -- CP-element group 879: 	882 
    -- CP-element group 879:  members (2) 
      -- CP-element group 879: 	 branch_block_stmt_223/merge_stmt_3063_PhiReqMerge
      -- CP-element group 879: 	 branch_block_stmt_223/merge_stmt_3063_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(879) <= OrReduce(zeropad3D_CP_676_elements(872) & zeropad3D_CP_676_elements(878));
    -- CP-element group 880:  transition  input  bypass 
    -- CP-element group 880: predecessors 
    -- CP-element group 880: 	879 
    -- CP-element group 880: successors 
    -- CP-element group 880: 	883 
    -- CP-element group 880:  members (1) 
      -- CP-element group 880: 	 branch_block_stmt_223/merge_stmt_3063_PhiAck/phi_stmt_3064_ack
      -- 
    phi_stmt_3064_ack_8853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 880_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3064_ack_0, ack => zeropad3D_CP_676_elements(880)); -- 
    -- CP-element group 881:  transition  input  bypass 
    -- CP-element group 881: predecessors 
    -- CP-element group 881: 	879 
    -- CP-element group 881: successors 
    -- CP-element group 881: 	883 
    -- CP-element group 881:  members (1) 
      -- CP-element group 881: 	 branch_block_stmt_223/merge_stmt_3063_PhiAck/phi_stmt_3071_ack
      -- 
    phi_stmt_3071_ack_8854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 881_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3071_ack_0, ack => zeropad3D_CP_676_elements(881)); -- 
    -- CP-element group 882:  transition  input  bypass 
    -- CP-element group 882: predecessors 
    -- CP-element group 882: 	879 
    -- CP-element group 882: successors 
    -- CP-element group 882: 	883 
    -- CP-element group 882:  members (1) 
      -- CP-element group 882: 	 branch_block_stmt_223/merge_stmt_3063_PhiAck/phi_stmt_3077_ack
      -- 
    phi_stmt_3077_ack_8855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 882_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3077_ack_0, ack => zeropad3D_CP_676_elements(882)); -- 
    -- CP-element group 883:  join  fork  transition  place  output  bypass 
    -- CP-element group 883: predecessors 
    -- CP-element group 883: 	880 
    -- CP-element group 883: 	881 
    -- CP-element group 883: 	882 
    -- CP-element group 883: successors 
    -- CP-element group 883: 	459 
    -- CP-element group 883: 	460 
    -- CP-element group 883:  members (10) 
      -- CP-element group 883: 	 branch_block_stmt_223/merge_stmt_3063__exit__
      -- CP-element group 883: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114__entry__
      -- CP-element group 883: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/$entry
      -- CP-element group 883: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_sample_start_
      -- CP-element group 883: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_update_start_
      -- CP-element group 883: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_Sample/$entry
      -- CP-element group 883: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_Sample/rr
      -- CP-element group 883: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_Update/$entry
      -- CP-element group 883: 	 branch_block_stmt_223/assign_stmt_3089_to_assign_stmt_3114/type_cast_3088_Update/cr
      -- CP-element group 883: 	 branch_block_stmt_223/merge_stmt_3063_PhiAck/$exit
      -- 
    rr_5442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(883), ack => type_cast_3088_inst_req_0); -- 
    cr_5447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(883), ack => type_cast_3088_inst_req_1); -- 
    zeropad3D_cp_element_group_883: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_883"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(880) & zeropad3D_CP_676_elements(881) & zeropad3D_CP_676_elements(882);
      gj_zeropad3D_cp_element_group_883 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(883), clk => clk, reset => reset); --
    end block;
    -- CP-element group 884:  merge  fork  transition  place  output  bypass 
    -- CP-element group 884: predecessors 
    -- CP-element group 884: 	462 
    -- CP-element group 884: 	466 
    -- CP-element group 884: successors 
    -- CP-element group 884: 	467 
    -- CP-element group 884: 	468 
    -- CP-element group 884: 	469 
    -- CP-element group 884: 	470 
    -- CP-element group 884: 	473 
    -- CP-element group 884: 	475 
    -- CP-element group 884: 	477 
    -- CP-element group 884: 	479 
    -- CP-element group 884:  members (33) 
      -- CP-element group 884: 	 branch_block_stmt_223/merge_stmt_3158__exit__
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214__entry__
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_sample_start_
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_update_start_
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_Sample/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_Sample/rr
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_Update/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3162_Update/cr
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_sample_start_
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_update_start_
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_Sample/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_Sample/rr
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_Update/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3167_Update/cr
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_update_start_
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_Update/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/type_cast_3201_Update/cr
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_update_start_
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_final_index_sum_regn_update_start
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_final_index_sum_regn_Update/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/array_obj_ref_3207_final_index_sum_regn_Update/req
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_complete/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/addr_of_3208_complete/req
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_update_start_
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Update/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Update/word_access_complete/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Update/word_access_complete/word_0/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/assign_stmt_3163_to_assign_stmt_3214/ptr_deref_3211_Update/word_access_complete/word_0/cr
      -- CP-element group 884: 	 branch_block_stmt_223/merge_stmt_3158_PhiReqMerge
      -- CP-element group 884: 	 branch_block_stmt_223/merge_stmt_3158_PhiAck/$entry
      -- CP-element group 884: 	 branch_block_stmt_223/merge_stmt_3158_PhiAck/$exit
      -- CP-element group 884: 	 branch_block_stmt_223/merge_stmt_3158_PhiAck/dummy
      -- 
    rr_5514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(884), ack => type_cast_3162_inst_req_0); -- 
    cr_5519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(884), ack => type_cast_3162_inst_req_1); -- 
    rr_5528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(884), ack => type_cast_3167_inst_req_0); -- 
    cr_5533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(884), ack => type_cast_3167_inst_req_1); -- 
    cr_5547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(884), ack => type_cast_3201_inst_req_1); -- 
    req_5578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(884), ack => array_obj_ref_3207_index_offset_req_1); -- 
    req_5593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(884), ack => addr_of_3208_final_reg_req_1); -- 
    cr_5643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(884), ack => ptr_deref_3211_store_0_req_1); -- 
    zeropad3D_CP_676_elements(884) <= OrReduce(zeropad3D_CP_676_elements(462) & zeropad3D_CP_676_elements(466));
    -- CP-element group 885:  merge  fork  transition  place  output  bypass 
    -- CP-element group 885: predecessors 
    -- CP-element group 885: 	480 
    -- CP-element group 885: 	500 
    -- CP-element group 885: successors 
    -- CP-element group 885: 	501 
    -- CP-element group 885: 	502 
    -- CP-element group 885:  members (13) 
      -- CP-element group 885: 	 branch_block_stmt_223/merge_stmt_3323__exit__
      -- CP-element group 885: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341__entry__
      -- CP-element group 885: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_sample_start_
      -- CP-element group 885: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_update_start_
      -- CP-element group 885: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_Sample/$entry
      -- CP-element group 885: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_Sample/rr
      -- CP-element group 885: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_Update/$entry
      -- CP-element group 885: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/type_cast_3327_Update/cr
      -- CP-element group 885: 	 branch_block_stmt_223/assign_stmt_3328_to_assign_stmt_3341/$entry
      -- CP-element group 885: 	 branch_block_stmt_223/merge_stmt_3323_PhiReqMerge
      -- CP-element group 885: 	 branch_block_stmt_223/merge_stmt_3323_PhiAck/$entry
      -- CP-element group 885: 	 branch_block_stmt_223/merge_stmt_3323_PhiAck/$exit
      -- CP-element group 885: 	 branch_block_stmt_223/merge_stmt_3323_PhiAck/dummy
      -- 
    rr_5892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(885), ack => type_cast_3327_inst_req_0); -- 
    cr_5897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(885), ack => type_cast_3327_inst_req_1); -- 
    zeropad3D_CP_676_elements(885) <= OrReduce(zeropad3D_CP_676_elements(480) & zeropad3D_CP_676_elements(500));
    -- CP-element group 886:  transition  input  bypass 
    -- CP-element group 886: predecessors 
    -- CP-element group 886: 	512 
    -- CP-element group 886: successors 
    -- CP-element group 886: 	888 
    -- CP-element group 886:  members (2) 
      -- CP-element group 886: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/SplitProtocol/Sample/$exit
      -- CP-element group 886: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/SplitProtocol/Sample/ra
      -- 
    ra_8945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 886_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3422_inst_ack_0, ack => zeropad3D_CP_676_elements(886)); -- 
    -- CP-element group 887:  transition  input  bypass 
    -- CP-element group 887: predecessors 
    -- CP-element group 887: 	512 
    -- CP-element group 887: successors 
    -- CP-element group 887: 	888 
    -- CP-element group 887:  members (2) 
      -- CP-element group 887: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/SplitProtocol/Update/$exit
      -- CP-element group 887: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/SplitProtocol/Update/ca
      -- 
    ca_8950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 887_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3422_inst_ack_1, ack => zeropad3D_CP_676_elements(887)); -- 
    -- CP-element group 888:  join  transition  output  bypass 
    -- CP-element group 888: predecessors 
    -- CP-element group 888: 	886 
    -- CP-element group 888: 	887 
    -- CP-element group 888: successors 
    -- CP-element group 888: 	893 
    -- CP-element group 888:  members (5) 
      -- CP-element group 888: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/$exit
      -- CP-element group 888: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/$exit
      -- CP-element group 888: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/$exit
      -- CP-element group 888: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3422/SplitProtocol/$exit
      -- CP-element group 888: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_req
      -- 
    phi_stmt_3419_req_8951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3419_req_8951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(888), ack => phi_stmt_3419_req_0); -- 
    zeropad3D_cp_element_group_888: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_888"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(886) & zeropad3D_CP_676_elements(887);
      gj_zeropad3D_cp_element_group_888 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(888), clk => clk, reset => reset); --
    end block;
    -- CP-element group 889:  transition  output  delay-element  bypass 
    -- CP-element group 889: predecessors 
    -- CP-element group 889: 	512 
    -- CP-element group 889: successors 
    -- CP-element group 889: 	893 
    -- CP-element group 889:  members (4) 
      -- CP-element group 889: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3406/$exit
      -- CP-element group 889: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/$exit
      -- CP-element group 889: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3410_konst_delay_trans
      -- CP-element group 889: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_req
      -- 
    phi_stmt_3406_req_8959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3406_req_8959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(889), ack => phi_stmt_3406_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(889) is a control-delay.
    cp_element_889_delay: control_delay_element  generic map(name => " 889_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(512), ack => zeropad3D_CP_676_elements(889), clk => clk, reset =>reset);
    -- CP-element group 890:  transition  input  bypass 
    -- CP-element group 890: predecessors 
    -- CP-element group 890: 	512 
    -- CP-element group 890: successors 
    -- CP-element group 890: 	892 
    -- CP-element group 890:  members (2) 
      -- CP-element group 890: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/SplitProtocol/Sample/$exit
      -- CP-element group 890: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/SplitProtocol/Sample/ra
      -- 
    ra_8976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 890_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3416_inst_ack_0, ack => zeropad3D_CP_676_elements(890)); -- 
    -- CP-element group 891:  transition  input  bypass 
    -- CP-element group 891: predecessors 
    -- CP-element group 891: 	512 
    -- CP-element group 891: successors 
    -- CP-element group 891: 	892 
    -- CP-element group 891:  members (2) 
      -- CP-element group 891: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/SplitProtocol/Update/$exit
      -- CP-element group 891: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/SplitProtocol/Update/ca
      -- 
    ca_8981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 891_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3416_inst_ack_1, ack => zeropad3D_CP_676_elements(891)); -- 
    -- CP-element group 892:  join  transition  output  bypass 
    -- CP-element group 892: predecessors 
    -- CP-element group 892: 	890 
    -- CP-element group 892: 	891 
    -- CP-element group 892: successors 
    -- CP-element group 892: 	893 
    -- CP-element group 892:  members (5) 
      -- CP-element group 892: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/$exit
      -- CP-element group 892: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/$exit
      -- CP-element group 892: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/$exit
      -- CP-element group 892: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3416/SplitProtocol/$exit
      -- CP-element group 892: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_req
      -- 
    phi_stmt_3413_req_8982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3413_req_8982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(892), ack => phi_stmt_3413_req_0); -- 
    zeropad3D_cp_element_group_892: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_892"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(890) & zeropad3D_CP_676_elements(891);
      gj_zeropad3D_cp_element_group_892 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(892), clk => clk, reset => reset); --
    end block;
    -- CP-element group 893:  join  transition  bypass 
    -- CP-element group 893: predecessors 
    -- CP-element group 893: 	888 
    -- CP-element group 893: 	889 
    -- CP-element group 893: 	892 
    -- CP-element group 893: successors 
    -- CP-element group 893: 	904 
    -- CP-element group 893:  members (1) 
      -- CP-element group 893: 	 branch_block_stmt_223/ifx_xelse1529_ifx_xend1565_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_893: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_893"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(888) & zeropad3D_CP_676_elements(889) & zeropad3D_CP_676_elements(892);
      gj_zeropad3D_cp_element_group_893 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(893), clk => clk, reset => reset); --
    end block;
    -- CP-element group 894:  transition  input  bypass 
    -- CP-element group 894: predecessors 
    -- CP-element group 894: 	503 
    -- CP-element group 894: successors 
    -- CP-element group 894: 	896 
    -- CP-element group 894:  members (2) 
      -- CP-element group 894: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/SplitProtocol/Sample/$exit
      -- CP-element group 894: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/SplitProtocol/Sample/ra
      -- 
    ra_9002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 894_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3424_inst_ack_0, ack => zeropad3D_CP_676_elements(894)); -- 
    -- CP-element group 895:  transition  input  bypass 
    -- CP-element group 895: predecessors 
    -- CP-element group 895: 	503 
    -- CP-element group 895: successors 
    -- CP-element group 895: 	896 
    -- CP-element group 895:  members (2) 
      -- CP-element group 895: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/SplitProtocol/Update/$exit
      -- CP-element group 895: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/SplitProtocol/Update/ca
      -- 
    ca_9007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 895_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3424_inst_ack_1, ack => zeropad3D_CP_676_elements(895)); -- 
    -- CP-element group 896:  join  transition  output  bypass 
    -- CP-element group 896: predecessors 
    -- CP-element group 896: 	894 
    -- CP-element group 896: 	895 
    -- CP-element group 896: successors 
    -- CP-element group 896: 	903 
    -- CP-element group 896:  members (5) 
      -- CP-element group 896: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/$exit
      -- CP-element group 896: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/$exit
      -- CP-element group 896: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/$exit
      -- CP-element group 896: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_sources/type_cast_3424/SplitProtocol/$exit
      -- CP-element group 896: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3419/phi_stmt_3419_req
      -- 
    phi_stmt_3419_req_9008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3419_req_9008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(896), ack => phi_stmt_3419_req_1); -- 
    zeropad3D_cp_element_group_896: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_896"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(894) & zeropad3D_CP_676_elements(895);
      gj_zeropad3D_cp_element_group_896 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(896), clk => clk, reset => reset); --
    end block;
    -- CP-element group 897:  transition  input  bypass 
    -- CP-element group 897: predecessors 
    -- CP-element group 897: 	503 
    -- CP-element group 897: successors 
    -- CP-element group 897: 	899 
    -- CP-element group 897:  members (2) 
      -- CP-element group 897: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/SplitProtocol/Sample/$exit
      -- CP-element group 897: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/SplitProtocol/Sample/ra
      -- 
    ra_9025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 897_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3412_inst_ack_0, ack => zeropad3D_CP_676_elements(897)); -- 
    -- CP-element group 898:  transition  input  bypass 
    -- CP-element group 898: predecessors 
    -- CP-element group 898: 	503 
    -- CP-element group 898: successors 
    -- CP-element group 898: 	899 
    -- CP-element group 898:  members (2) 
      -- CP-element group 898: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/SplitProtocol/Update/$exit
      -- CP-element group 898: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/SplitProtocol/Update/ca
      -- 
    ca_9030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 898_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3412_inst_ack_1, ack => zeropad3D_CP_676_elements(898)); -- 
    -- CP-element group 899:  join  transition  output  bypass 
    -- CP-element group 899: predecessors 
    -- CP-element group 899: 	897 
    -- CP-element group 899: 	898 
    -- CP-element group 899: successors 
    -- CP-element group 899: 	903 
    -- CP-element group 899:  members (5) 
      -- CP-element group 899: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/$exit
      -- CP-element group 899: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/$exit
      -- CP-element group 899: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/$exit
      -- CP-element group 899: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_sources/type_cast_3412/SplitProtocol/$exit
      -- CP-element group 899: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3406/phi_stmt_3406_req
      -- 
    phi_stmt_3406_req_9031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3406_req_9031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(899), ack => phi_stmt_3406_req_1); -- 
    zeropad3D_cp_element_group_899: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_899"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(897) & zeropad3D_CP_676_elements(898);
      gj_zeropad3D_cp_element_group_899 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(899), clk => clk, reset => reset); --
    end block;
    -- CP-element group 900:  transition  input  bypass 
    -- CP-element group 900: predecessors 
    -- CP-element group 900: 	503 
    -- CP-element group 900: successors 
    -- CP-element group 900: 	902 
    -- CP-element group 900:  members (2) 
      -- CP-element group 900: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/SplitProtocol/Sample/$exit
      -- CP-element group 900: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/SplitProtocol/Sample/ra
      -- 
    ra_9048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 900_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3418_inst_ack_0, ack => zeropad3D_CP_676_elements(900)); -- 
    -- CP-element group 901:  transition  input  bypass 
    -- CP-element group 901: predecessors 
    -- CP-element group 901: 	503 
    -- CP-element group 901: successors 
    -- CP-element group 901: 	902 
    -- CP-element group 901:  members (2) 
      -- CP-element group 901: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/SplitProtocol/Update/$exit
      -- CP-element group 901: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/SplitProtocol/Update/ca
      -- 
    ca_9053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 901_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3418_inst_ack_1, ack => zeropad3D_CP_676_elements(901)); -- 
    -- CP-element group 902:  join  transition  output  bypass 
    -- CP-element group 902: predecessors 
    -- CP-element group 902: 	900 
    -- CP-element group 902: 	901 
    -- CP-element group 902: successors 
    -- CP-element group 902: 	903 
    -- CP-element group 902:  members (5) 
      -- CP-element group 902: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/$exit
      -- CP-element group 902: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/$exit
      -- CP-element group 902: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/$exit
      -- CP-element group 902: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_sources/type_cast_3418/SplitProtocol/$exit
      -- CP-element group 902: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/phi_stmt_3413/phi_stmt_3413_req
      -- 
    phi_stmt_3413_req_9054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3413_req_9054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(902), ack => phi_stmt_3413_req_1); -- 
    zeropad3D_cp_element_group_902: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_902"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(900) & zeropad3D_CP_676_elements(901);
      gj_zeropad3D_cp_element_group_902 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(902), clk => clk, reset => reset); --
    end block;
    -- CP-element group 903:  join  transition  bypass 
    -- CP-element group 903: predecessors 
    -- CP-element group 903: 	896 
    -- CP-element group 903: 	899 
    -- CP-element group 903: 	902 
    -- CP-element group 903: successors 
    -- CP-element group 903: 	904 
    -- CP-element group 903:  members (1) 
      -- CP-element group 903: 	 branch_block_stmt_223/ifx_xthen1524_ifx_xend1565_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_903: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_903"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(896) & zeropad3D_CP_676_elements(899) & zeropad3D_CP_676_elements(902);
      gj_zeropad3D_cp_element_group_903 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(903), clk => clk, reset => reset); --
    end block;
    -- CP-element group 904:  merge  fork  transition  place  bypass 
    -- CP-element group 904: predecessors 
    -- CP-element group 904: 	893 
    -- CP-element group 904: 	903 
    -- CP-element group 904: successors 
    -- CP-element group 904: 	905 
    -- CP-element group 904: 	906 
    -- CP-element group 904: 	907 
    -- CP-element group 904:  members (2) 
      -- CP-element group 904: 	 branch_block_stmt_223/merge_stmt_3405_PhiReqMerge
      -- CP-element group 904: 	 branch_block_stmt_223/merge_stmt_3405_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(904) <= OrReduce(zeropad3D_CP_676_elements(893) & zeropad3D_CP_676_elements(903));
    -- CP-element group 905:  transition  input  bypass 
    -- CP-element group 905: predecessors 
    -- CP-element group 905: 	904 
    -- CP-element group 905: successors 
    -- CP-element group 905: 	908 
    -- CP-element group 905:  members (1) 
      -- CP-element group 905: 	 branch_block_stmt_223/merge_stmt_3405_PhiAck/phi_stmt_3406_ack
      -- 
    phi_stmt_3406_ack_9059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 905_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3406_ack_0, ack => zeropad3D_CP_676_elements(905)); -- 
    -- CP-element group 906:  transition  input  bypass 
    -- CP-element group 906: predecessors 
    -- CP-element group 906: 	904 
    -- CP-element group 906: successors 
    -- CP-element group 906: 	908 
    -- CP-element group 906:  members (1) 
      -- CP-element group 906: 	 branch_block_stmt_223/merge_stmt_3405_PhiAck/phi_stmt_3413_ack
      -- 
    phi_stmt_3413_ack_9060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 906_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3413_ack_0, ack => zeropad3D_CP_676_elements(906)); -- 
    -- CP-element group 907:  transition  input  bypass 
    -- CP-element group 907: predecessors 
    -- CP-element group 907: 	904 
    -- CP-element group 907: successors 
    -- CP-element group 907: 	908 
    -- CP-element group 907:  members (1) 
      -- CP-element group 907: 	 branch_block_stmt_223/merge_stmt_3405_PhiAck/phi_stmt_3419_ack
      -- 
    phi_stmt_3419_ack_9061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 907_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3419_ack_0, ack => zeropad3D_CP_676_elements(907)); -- 
    -- CP-element group 908:  join  transition  bypass 
    -- CP-element group 908: predecessors 
    -- CP-element group 908: 	905 
    -- CP-element group 908: 	906 
    -- CP-element group 908: 	907 
    -- CP-element group 908: successors 
    -- CP-element group 908: 	7 
    -- CP-element group 908:  members (1) 
      -- CP-element group 908: 	 branch_block_stmt_223/merge_stmt_3405_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_908: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_908"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(905) & zeropad3D_CP_676_elements(906) & zeropad3D_CP_676_elements(907);
      gj_zeropad3D_cp_element_group_908 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(908), clk => clk, reset => reset); --
    end block;
    -- CP-element group 909:  transition  input  bypass 
    -- CP-element group 909: predecessors 
    -- CP-element group 909: 	8 
    -- CP-element group 909: successors 
    -- CP-element group 909: 	911 
    -- CP-element group 909:  members (2) 
      -- CP-element group 909: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/SplitProtocol/Sample/$exit
      -- CP-element group 909: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/SplitProtocol/Sample/ra
      -- 
    ra_9089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 909_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3481_inst_ack_0, ack => zeropad3D_CP_676_elements(909)); -- 
    -- CP-element group 910:  transition  input  bypass 
    -- CP-element group 910: predecessors 
    -- CP-element group 910: 	8 
    -- CP-element group 910: successors 
    -- CP-element group 910: 	911 
    -- CP-element group 910:  members (2) 
      -- CP-element group 910: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/SplitProtocol/Update/$exit
      -- CP-element group 910: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/SplitProtocol/Update/ca
      -- 
    ca_9094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 910_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3481_inst_ack_1, ack => zeropad3D_CP_676_elements(910)); -- 
    -- CP-element group 911:  join  transition  output  bypass 
    -- CP-element group 911: predecessors 
    -- CP-element group 911: 	909 
    -- CP-element group 911: 	910 
    -- CP-element group 911: successors 
    -- CP-element group 911: 	918 
    -- CP-element group 911:  members (5) 
      -- CP-element group 911: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/$exit
      -- CP-element group 911: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/$exit
      -- CP-element group 911: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/$exit
      -- CP-element group 911: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3481/SplitProtocol/$exit
      -- CP-element group 911: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_req
      -- 
    phi_stmt_3475_req_9095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3475_req_9095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(911), ack => phi_stmt_3475_req_1); -- 
    zeropad3D_cp_element_group_911: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_911"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(909) & zeropad3D_CP_676_elements(910);
      gj_zeropad3D_cp_element_group_911 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(911), clk => clk, reset => reset); --
    end block;
    -- CP-element group 912:  transition  input  bypass 
    -- CP-element group 912: predecessors 
    -- CP-element group 912: 	8 
    -- CP-element group 912: successors 
    -- CP-element group 912: 	914 
    -- CP-element group 912:  members (2) 
      -- CP-element group 912: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/SplitProtocol/Sample/$exit
      -- CP-element group 912: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/SplitProtocol/Sample/ra
      -- 
    ra_9112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 912_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3487_inst_ack_0, ack => zeropad3D_CP_676_elements(912)); -- 
    -- CP-element group 913:  transition  input  bypass 
    -- CP-element group 913: predecessors 
    -- CP-element group 913: 	8 
    -- CP-element group 913: successors 
    -- CP-element group 913: 	914 
    -- CP-element group 913:  members (2) 
      -- CP-element group 913: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/SplitProtocol/Update/$exit
      -- CP-element group 913: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/SplitProtocol/Update/ca
      -- 
    ca_9117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 913_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3487_inst_ack_1, ack => zeropad3D_CP_676_elements(913)); -- 
    -- CP-element group 914:  join  transition  output  bypass 
    -- CP-element group 914: predecessors 
    -- CP-element group 914: 	912 
    -- CP-element group 914: 	913 
    -- CP-element group 914: successors 
    -- CP-element group 914: 	918 
    -- CP-element group 914:  members (5) 
      -- CP-element group 914: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/$exit
      -- CP-element group 914: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/$exit
      -- CP-element group 914: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/$exit
      -- CP-element group 914: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3487/SplitProtocol/$exit
      -- CP-element group 914: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_req
      -- 
    phi_stmt_3482_req_9118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3482_req_9118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(914), ack => phi_stmt_3482_req_1); -- 
    zeropad3D_cp_element_group_914: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_914"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(912) & zeropad3D_CP_676_elements(913);
      gj_zeropad3D_cp_element_group_914 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(914), clk => clk, reset => reset); --
    end block;
    -- CP-element group 915:  transition  input  bypass 
    -- CP-element group 915: predecessors 
    -- CP-element group 915: 	8 
    -- CP-element group 915: successors 
    -- CP-element group 915: 	917 
    -- CP-element group 915:  members (2) 
      -- CP-element group 915: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/SplitProtocol/Sample/$exit
      -- CP-element group 915: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/SplitProtocol/Sample/ra
      -- 
    ra_9135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 915_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3493_inst_ack_0, ack => zeropad3D_CP_676_elements(915)); -- 
    -- CP-element group 916:  transition  input  bypass 
    -- CP-element group 916: predecessors 
    -- CP-element group 916: 	8 
    -- CP-element group 916: successors 
    -- CP-element group 916: 	917 
    -- CP-element group 916:  members (2) 
      -- CP-element group 916: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/SplitProtocol/Update/$exit
      -- CP-element group 916: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/SplitProtocol/Update/ca
      -- 
    ca_9140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 916_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3493_inst_ack_1, ack => zeropad3D_CP_676_elements(916)); -- 
    -- CP-element group 917:  join  transition  output  bypass 
    -- CP-element group 917: predecessors 
    -- CP-element group 917: 	915 
    -- CP-element group 917: 	916 
    -- CP-element group 917: successors 
    -- CP-element group 917: 	918 
    -- CP-element group 917:  members (5) 
      -- CP-element group 917: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/$exit
      -- CP-element group 917: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/$exit
      -- CP-element group 917: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/$exit
      -- CP-element group 917: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3493/SplitProtocol/$exit
      -- CP-element group 917: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_req
      -- 
    phi_stmt_3488_req_9141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3488_req_9141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(917), ack => phi_stmt_3488_req_1); -- 
    zeropad3D_cp_element_group_917: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_917"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(915) & zeropad3D_CP_676_elements(916);
      gj_zeropad3D_cp_element_group_917 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(917), clk => clk, reset => reset); --
    end block;
    -- CP-element group 918:  join  transition  bypass 
    -- CP-element group 918: predecessors 
    -- CP-element group 918: 	911 
    -- CP-element group 918: 	914 
    -- CP-element group 918: 	917 
    -- CP-element group 918: successors 
    -- CP-element group 918: 	927 
    -- CP-element group 918:  members (1) 
      -- CP-element group 918: 	 branch_block_stmt_223/ifx_xend1784_whilex_xbody1631_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_918: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_918"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(911) & zeropad3D_CP_676_elements(914) & zeropad3D_CP_676_elements(917);
      gj_zeropad3D_cp_element_group_918 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(918), clk => clk, reset => reset); --
    end block;
    -- CP-element group 919:  transition  output  delay-element  bypass 
    -- CP-element group 919: predecessors 
    -- CP-element group 919: 	516 
    -- CP-element group 919: successors 
    -- CP-element group 919: 	926 
    -- CP-element group 919:  members (4) 
      -- CP-element group 919: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3475/$exit
      -- CP-element group 919: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/$exit
      -- CP-element group 919: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_sources/type_cast_3479_konst_delay_trans
      -- CP-element group 919: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3475/phi_stmt_3475_req
      -- 
    phi_stmt_3475_req_9152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3475_req_9152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(919), ack => phi_stmt_3475_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(919) is a control-delay.
    cp_element_919_delay: control_delay_element  generic map(name => " 919_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(516), ack => zeropad3D_CP_676_elements(919), clk => clk, reset =>reset);
    -- CP-element group 920:  transition  input  bypass 
    -- CP-element group 920: predecessors 
    -- CP-element group 920: 	516 
    -- CP-element group 920: successors 
    -- CP-element group 920: 	922 
    -- CP-element group 920:  members (2) 
      -- CP-element group 920: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/SplitProtocol/Sample/$exit
      -- CP-element group 920: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/SplitProtocol/Sample/ra
      -- 
    ra_9169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 920_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3485_inst_ack_0, ack => zeropad3D_CP_676_elements(920)); -- 
    -- CP-element group 921:  transition  input  bypass 
    -- CP-element group 921: predecessors 
    -- CP-element group 921: 	516 
    -- CP-element group 921: successors 
    -- CP-element group 921: 	922 
    -- CP-element group 921:  members (2) 
      -- CP-element group 921: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/SplitProtocol/Update/$exit
      -- CP-element group 921: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/SplitProtocol/Update/ca
      -- 
    ca_9174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 921_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3485_inst_ack_1, ack => zeropad3D_CP_676_elements(921)); -- 
    -- CP-element group 922:  join  transition  output  bypass 
    -- CP-element group 922: predecessors 
    -- CP-element group 922: 	920 
    -- CP-element group 922: 	921 
    -- CP-element group 922: successors 
    -- CP-element group 922: 	926 
    -- CP-element group 922:  members (5) 
      -- CP-element group 922: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/$exit
      -- CP-element group 922: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/$exit
      -- CP-element group 922: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/$exit
      -- CP-element group 922: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_sources/type_cast_3485/SplitProtocol/$exit
      -- CP-element group 922: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3482/phi_stmt_3482_req
      -- 
    phi_stmt_3482_req_9175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3482_req_9175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(922), ack => phi_stmt_3482_req_0); -- 
    zeropad3D_cp_element_group_922: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_922"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(920) & zeropad3D_CP_676_elements(921);
      gj_zeropad3D_cp_element_group_922 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(922), clk => clk, reset => reset); --
    end block;
    -- CP-element group 923:  transition  input  bypass 
    -- CP-element group 923: predecessors 
    -- CP-element group 923: 	516 
    -- CP-element group 923: successors 
    -- CP-element group 923: 	925 
    -- CP-element group 923:  members (2) 
      -- CP-element group 923: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/SplitProtocol/Sample/$exit
      -- CP-element group 923: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/SplitProtocol/Sample/ra
      -- 
    ra_9192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 923_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3491_inst_ack_0, ack => zeropad3D_CP_676_elements(923)); -- 
    -- CP-element group 924:  transition  input  bypass 
    -- CP-element group 924: predecessors 
    -- CP-element group 924: 	516 
    -- CP-element group 924: successors 
    -- CP-element group 924: 	925 
    -- CP-element group 924:  members (2) 
      -- CP-element group 924: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/SplitProtocol/Update/$exit
      -- CP-element group 924: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/SplitProtocol/Update/ca
      -- 
    ca_9197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 924_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3491_inst_ack_1, ack => zeropad3D_CP_676_elements(924)); -- 
    -- CP-element group 925:  join  transition  output  bypass 
    -- CP-element group 925: predecessors 
    -- CP-element group 925: 	923 
    -- CP-element group 925: 	924 
    -- CP-element group 925: successors 
    -- CP-element group 925: 	926 
    -- CP-element group 925:  members (5) 
      -- CP-element group 925: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/$exit
      -- CP-element group 925: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/$exit
      -- CP-element group 925: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/$exit
      -- CP-element group 925: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_sources/type_cast_3491/SplitProtocol/$exit
      -- CP-element group 925: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/phi_stmt_3488/phi_stmt_3488_req
      -- 
    phi_stmt_3488_req_9198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3488_req_9198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(925), ack => phi_stmt_3488_req_0); -- 
    zeropad3D_cp_element_group_925: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_925"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(923) & zeropad3D_CP_676_elements(924);
      gj_zeropad3D_cp_element_group_925 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(925), clk => clk, reset => reset); --
    end block;
    -- CP-element group 926:  join  transition  bypass 
    -- CP-element group 926: predecessors 
    -- CP-element group 926: 	919 
    -- CP-element group 926: 	922 
    -- CP-element group 926: 	925 
    -- CP-element group 926: successors 
    -- CP-element group 926: 	927 
    -- CP-element group 926:  members (1) 
      -- CP-element group 926: 	 branch_block_stmt_223/whilex_xend1566_whilex_xbody1631_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_926: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_926"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(919) & zeropad3D_CP_676_elements(922) & zeropad3D_CP_676_elements(925);
      gj_zeropad3D_cp_element_group_926 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(926), clk => clk, reset => reset); --
    end block;
    -- CP-element group 927:  merge  fork  transition  place  bypass 
    -- CP-element group 927: predecessors 
    -- CP-element group 927: 	918 
    -- CP-element group 927: 	926 
    -- CP-element group 927: successors 
    -- CP-element group 927: 	928 
    -- CP-element group 927: 	929 
    -- CP-element group 927: 	930 
    -- CP-element group 927:  members (2) 
      -- CP-element group 927: 	 branch_block_stmt_223/merge_stmt_3474_PhiReqMerge
      -- CP-element group 927: 	 branch_block_stmt_223/merge_stmt_3474_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(927) <= OrReduce(zeropad3D_CP_676_elements(918) & zeropad3D_CP_676_elements(926));
    -- CP-element group 928:  transition  input  bypass 
    -- CP-element group 928: predecessors 
    -- CP-element group 928: 	927 
    -- CP-element group 928: successors 
    -- CP-element group 928: 	931 
    -- CP-element group 928:  members (1) 
      -- CP-element group 928: 	 branch_block_stmt_223/merge_stmt_3474_PhiAck/phi_stmt_3475_ack
      -- 
    phi_stmt_3475_ack_9203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 928_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3475_ack_0, ack => zeropad3D_CP_676_elements(928)); -- 
    -- CP-element group 929:  transition  input  bypass 
    -- CP-element group 929: predecessors 
    -- CP-element group 929: 	927 
    -- CP-element group 929: successors 
    -- CP-element group 929: 	931 
    -- CP-element group 929:  members (1) 
      -- CP-element group 929: 	 branch_block_stmt_223/merge_stmt_3474_PhiAck/phi_stmt_3482_ack
      -- 
    phi_stmt_3482_ack_9204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 929_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3482_ack_0, ack => zeropad3D_CP_676_elements(929)); -- 
    -- CP-element group 930:  transition  input  bypass 
    -- CP-element group 930: predecessors 
    -- CP-element group 930: 	927 
    -- CP-element group 930: successors 
    -- CP-element group 930: 	931 
    -- CP-element group 930:  members (1) 
      -- CP-element group 930: 	 branch_block_stmt_223/merge_stmt_3474_PhiAck/phi_stmt_3488_ack
      -- 
    phi_stmt_3488_ack_9205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 930_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3488_ack_0, ack => zeropad3D_CP_676_elements(930)); -- 
    -- CP-element group 931:  join  fork  transition  place  output  bypass 
    -- CP-element group 931: predecessors 
    -- CP-element group 931: 	928 
    -- CP-element group 931: 	929 
    -- CP-element group 931: 	930 
    -- CP-element group 931: successors 
    -- CP-element group 931: 	517 
    -- CP-element group 931: 	518 
    -- CP-element group 931:  members (10) 
      -- CP-element group 931: 	 branch_block_stmt_223/merge_stmt_3474__exit__
      -- CP-element group 931: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524__entry__
      -- CP-element group 931: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_Sample/$entry
      -- CP-element group 931: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_Sample/rr
      -- CP-element group 931: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_Update/$entry
      -- CP-element group 931: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_Update/cr
      -- CP-element group 931: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_update_start_
      -- CP-element group 931: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/type_cast_3498_sample_start_
      -- CP-element group 931: 	 branch_block_stmt_223/assign_stmt_3499_to_assign_stmt_3524/$entry
      -- CP-element group 931: 	 branch_block_stmt_223/merge_stmt_3474_PhiAck/$exit
      -- 
    rr_6045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(931), ack => type_cast_3498_inst_req_0); -- 
    cr_6050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(931), ack => type_cast_3498_inst_req_1); -- 
    zeropad3D_cp_element_group_931: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_931"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(928) & zeropad3D_CP_676_elements(929) & zeropad3D_CP_676_elements(930);
      gj_zeropad3D_cp_element_group_931 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(931), clk => clk, reset => reset); --
    end block;
    -- CP-element group 932:  merge  fork  transition  place  output  bypass 
    -- CP-element group 932: predecessors 
    -- CP-element group 932: 	520 
    -- CP-element group 932: 	524 
    -- CP-element group 932: successors 
    -- CP-element group 932: 	525 
    -- CP-element group 932: 	526 
    -- CP-element group 932: 	527 
    -- CP-element group 932: 	528 
    -- CP-element group 932: 	531 
    -- CP-element group 932: 	533 
    -- CP-element group 932: 	535 
    -- CP-element group 932: 	537 
    -- CP-element group 932:  members (33) 
      -- CP-element group 932: 	 branch_block_stmt_223/merge_stmt_3568__exit__
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624__entry__
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_sample_start_
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_update_start_
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_update_start_
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_Sample/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_update_start_
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_Update/cr
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_Update/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_sample_start_
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3611_update_start_
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_Update/cr
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_Update/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_Update/cr
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_Sample/rr
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3577_Sample/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_Update/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/type_cast_3572_Sample/rr
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_final_index_sum_regn_update_start
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_final_index_sum_regn_Update/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/array_obj_ref_3617_final_index_sum_regn_Update/req
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_complete/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/addr_of_3618_complete/req
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_update_start_
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Update/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Update/word_access_complete/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Update/word_access_complete/word_0/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/assign_stmt_3573_to_assign_stmt_3624/ptr_deref_3621_Update/word_access_complete/word_0/cr
      -- CP-element group 932: 	 branch_block_stmt_223/merge_stmt_3568_PhiReqMerge
      -- CP-element group 932: 	 branch_block_stmt_223/merge_stmt_3568_PhiAck/$entry
      -- CP-element group 932: 	 branch_block_stmt_223/merge_stmt_3568_PhiAck/$exit
      -- CP-element group 932: 	 branch_block_stmt_223/merge_stmt_3568_PhiAck/dummy
      -- 
    cr_6150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(932), ack => type_cast_3611_inst_req_1); -- 
    cr_6136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(932), ack => type_cast_3577_inst_req_1); -- 
    cr_6122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(932), ack => type_cast_3572_inst_req_1); -- 
    rr_6131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(932), ack => type_cast_3577_inst_req_0); -- 
    rr_6117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(932), ack => type_cast_3572_inst_req_0); -- 
    req_6181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(932), ack => array_obj_ref_3617_index_offset_req_1); -- 
    req_6196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(932), ack => addr_of_3618_final_reg_req_1); -- 
    cr_6246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(932), ack => ptr_deref_3621_store_0_req_1); -- 
    zeropad3D_CP_676_elements(932) <= OrReduce(zeropad3D_CP_676_elements(520) & zeropad3D_CP_676_elements(524));
    -- CP-element group 933:  merge  fork  transition  place  output  bypass 
    -- CP-element group 933: predecessors 
    -- CP-element group 933: 	538 
    -- CP-element group 933: 	558 
    -- CP-element group 933: successors 
    -- CP-element group 933: 	559 
    -- CP-element group 933: 	560 
    -- CP-element group 933:  members (13) 
      -- CP-element group 933: 	 branch_block_stmt_223/merge_stmt_3733__exit__
      -- CP-element group 933: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751__entry__
      -- CP-element group 933: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/$entry
      -- CP-element group 933: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_sample_start_
      -- CP-element group 933: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_update_start_
      -- CP-element group 933: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_Sample/$entry
      -- CP-element group 933: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_Sample/rr
      -- CP-element group 933: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_Update/$entry
      -- CP-element group 933: 	 branch_block_stmt_223/assign_stmt_3738_to_assign_stmt_3751/type_cast_3737_Update/cr
      -- CP-element group 933: 	 branch_block_stmt_223/merge_stmt_3733_PhiReqMerge
      -- CP-element group 933: 	 branch_block_stmt_223/merge_stmt_3733_PhiAck/$entry
      -- CP-element group 933: 	 branch_block_stmt_223/merge_stmt_3733_PhiAck/$exit
      -- CP-element group 933: 	 branch_block_stmt_223/merge_stmt_3733_PhiAck/dummy
      -- 
    rr_6495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(933), ack => type_cast_3737_inst_req_0); -- 
    cr_6500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(933), ack => type_cast_3737_inst_req_1); -- 
    zeropad3D_CP_676_elements(933) <= OrReduce(zeropad3D_CP_676_elements(538) & zeropad3D_CP_676_elements(558));
    -- CP-element group 934:  transition  output  delay-element  bypass 
    -- CP-element group 934: predecessors 
    -- CP-element group 934: 	570 
    -- CP-element group 934: successors 
    -- CP-element group 934: 	941 
    -- CP-element group 934:  members (4) 
      -- CP-element group 934: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3815/$exit
      -- CP-element group 934: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/$exit
      -- CP-element group 934: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3819_konst_delay_trans
      -- CP-element group 934: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_req
      -- 
    phi_stmt_3815_req_9286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3815_req_9286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(934), ack => phi_stmt_3815_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(934) is a control-delay.
    cp_element_934_delay: control_delay_element  generic map(name => " 934_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(570), ack => zeropad3D_CP_676_elements(934), clk => clk, reset =>reset);
    -- CP-element group 935:  transition  input  bypass 
    -- CP-element group 935: predecessors 
    -- CP-element group 935: 	570 
    -- CP-element group 935: successors 
    -- CP-element group 935: 	937 
    -- CP-element group 935:  members (2) 
      -- CP-element group 935: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/SplitProtocol/Sample/$exit
      -- CP-element group 935: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/SplitProtocol/Sample/ra
      -- 
    ra_9303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 935_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3827_inst_ack_0, ack => zeropad3D_CP_676_elements(935)); -- 
    -- CP-element group 936:  transition  input  bypass 
    -- CP-element group 936: predecessors 
    -- CP-element group 936: 	570 
    -- CP-element group 936: successors 
    -- CP-element group 936: 	937 
    -- CP-element group 936:  members (2) 
      -- CP-element group 936: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/SplitProtocol/Update/$exit
      -- CP-element group 936: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/SplitProtocol/Update/ca
      -- 
    ca_9308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 936_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3827_inst_ack_1, ack => zeropad3D_CP_676_elements(936)); -- 
    -- CP-element group 937:  join  transition  output  bypass 
    -- CP-element group 937: predecessors 
    -- CP-element group 937: 	935 
    -- CP-element group 937: 	936 
    -- CP-element group 937: successors 
    -- CP-element group 937: 	941 
    -- CP-element group 937:  members (5) 
      -- CP-element group 937: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/$exit
      -- CP-element group 937: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/$exit
      -- CP-element group 937: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/$exit
      -- CP-element group 937: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3827/SplitProtocol/$exit
      -- CP-element group 937: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_req
      -- 
    phi_stmt_3822_req_9309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3822_req_9309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(937), ack => phi_stmt_3822_req_1); -- 
    zeropad3D_cp_element_group_937: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_937"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(935) & zeropad3D_CP_676_elements(936);
      gj_zeropad3D_cp_element_group_937 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(937), clk => clk, reset => reset); --
    end block;
    -- CP-element group 938:  transition  input  bypass 
    -- CP-element group 938: predecessors 
    -- CP-element group 938: 	570 
    -- CP-element group 938: successors 
    -- CP-element group 938: 	940 
    -- CP-element group 938:  members (2) 
      -- CP-element group 938: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/SplitProtocol/Sample/$exit
      -- CP-element group 938: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/SplitProtocol/Sample/ra
      -- 
    ra_9326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 938_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3831_inst_ack_0, ack => zeropad3D_CP_676_elements(938)); -- 
    -- CP-element group 939:  transition  input  bypass 
    -- CP-element group 939: predecessors 
    -- CP-element group 939: 	570 
    -- CP-element group 939: successors 
    -- CP-element group 939: 	940 
    -- CP-element group 939:  members (2) 
      -- CP-element group 939: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/SplitProtocol/Update/$exit
      -- CP-element group 939: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/SplitProtocol/Update/ca
      -- 
    ca_9331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 939_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3831_inst_ack_1, ack => zeropad3D_CP_676_elements(939)); -- 
    -- CP-element group 940:  join  transition  output  bypass 
    -- CP-element group 940: predecessors 
    -- CP-element group 940: 	938 
    -- CP-element group 940: 	939 
    -- CP-element group 940: successors 
    -- CP-element group 940: 	941 
    -- CP-element group 940:  members (5) 
      -- CP-element group 940: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/$exit
      -- CP-element group 940: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/$exit
      -- CP-element group 940: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/$exit
      -- CP-element group 940: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3831/SplitProtocol/$exit
      -- CP-element group 940: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_req
      -- 
    phi_stmt_3828_req_9332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3828_req_9332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(940), ack => phi_stmt_3828_req_0); -- 
    zeropad3D_cp_element_group_940: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_940"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(938) & zeropad3D_CP_676_elements(939);
      gj_zeropad3D_cp_element_group_940 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(940), clk => clk, reset => reset); --
    end block;
    -- CP-element group 941:  join  transition  bypass 
    -- CP-element group 941: predecessors 
    -- CP-element group 941: 	934 
    -- CP-element group 941: 	937 
    -- CP-element group 941: 	940 
    -- CP-element group 941: successors 
    -- CP-element group 941: 	952 
    -- CP-element group 941:  members (1) 
      -- CP-element group 941: 	 branch_block_stmt_223/ifx_xelse1749_ifx_xend1784_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_941: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_941"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(934) & zeropad3D_CP_676_elements(937) & zeropad3D_CP_676_elements(940);
      gj_zeropad3D_cp_element_group_941 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(941), clk => clk, reset => reset); --
    end block;
    -- CP-element group 942:  transition  input  bypass 
    -- CP-element group 942: predecessors 
    -- CP-element group 942: 	561 
    -- CP-element group 942: successors 
    -- CP-element group 942: 	944 
    -- CP-element group 942:  members (2) 
      -- CP-element group 942: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/SplitProtocol/Sample/$exit
      -- CP-element group 942: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/SplitProtocol/Sample/ra
      -- 
    ra_9352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 942_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3821_inst_ack_0, ack => zeropad3D_CP_676_elements(942)); -- 
    -- CP-element group 943:  transition  input  bypass 
    -- CP-element group 943: predecessors 
    -- CP-element group 943: 	561 
    -- CP-element group 943: successors 
    -- CP-element group 943: 	944 
    -- CP-element group 943:  members (2) 
      -- CP-element group 943: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/SplitProtocol/Update/$exit
      -- CP-element group 943: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/SplitProtocol/Update/ca
      -- 
    ca_9357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 943_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3821_inst_ack_1, ack => zeropad3D_CP_676_elements(943)); -- 
    -- CP-element group 944:  join  transition  output  bypass 
    -- CP-element group 944: predecessors 
    -- CP-element group 944: 	942 
    -- CP-element group 944: 	943 
    -- CP-element group 944: successors 
    -- CP-element group 944: 	951 
    -- CP-element group 944:  members (5) 
      -- CP-element group 944: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/$exit
      -- CP-element group 944: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/$exit
      -- CP-element group 944: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/$exit
      -- CP-element group 944: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_sources/type_cast_3821/SplitProtocol/$exit
      -- CP-element group 944: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3815/phi_stmt_3815_req
      -- 
    phi_stmt_3815_req_9358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3815_req_9358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(944), ack => phi_stmt_3815_req_1); -- 
    zeropad3D_cp_element_group_944: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_944"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(942) & zeropad3D_CP_676_elements(943);
      gj_zeropad3D_cp_element_group_944 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(944), clk => clk, reset => reset); --
    end block;
    -- CP-element group 945:  transition  input  bypass 
    -- CP-element group 945: predecessors 
    -- CP-element group 945: 	561 
    -- CP-element group 945: successors 
    -- CP-element group 945: 	947 
    -- CP-element group 945:  members (2) 
      -- CP-element group 945: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/SplitProtocol/Sample/$exit
      -- CP-element group 945: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/SplitProtocol/Sample/ra
      -- 
    ra_9375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 945_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3825_inst_ack_0, ack => zeropad3D_CP_676_elements(945)); -- 
    -- CP-element group 946:  transition  input  bypass 
    -- CP-element group 946: predecessors 
    -- CP-element group 946: 	561 
    -- CP-element group 946: successors 
    -- CP-element group 946: 	947 
    -- CP-element group 946:  members (2) 
      -- CP-element group 946: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/SplitProtocol/Update/$exit
      -- CP-element group 946: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/SplitProtocol/Update/ca
      -- 
    ca_9380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 946_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3825_inst_ack_1, ack => zeropad3D_CP_676_elements(946)); -- 
    -- CP-element group 947:  join  transition  output  bypass 
    -- CP-element group 947: predecessors 
    -- CP-element group 947: 	945 
    -- CP-element group 947: 	946 
    -- CP-element group 947: successors 
    -- CP-element group 947: 	951 
    -- CP-element group 947:  members (5) 
      -- CP-element group 947: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/$exit
      -- CP-element group 947: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/$exit
      -- CP-element group 947: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/$exit
      -- CP-element group 947: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_sources/type_cast_3825/SplitProtocol/$exit
      -- CP-element group 947: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3822/phi_stmt_3822_req
      -- 
    phi_stmt_3822_req_9381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3822_req_9381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(947), ack => phi_stmt_3822_req_0); -- 
    zeropad3D_cp_element_group_947: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_947"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(945) & zeropad3D_CP_676_elements(946);
      gj_zeropad3D_cp_element_group_947 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(947), clk => clk, reset => reset); --
    end block;
    -- CP-element group 948:  transition  input  bypass 
    -- CP-element group 948: predecessors 
    -- CP-element group 948: 	561 
    -- CP-element group 948: successors 
    -- CP-element group 948: 	950 
    -- CP-element group 948:  members (2) 
      -- CP-element group 948: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/SplitProtocol/Sample/$exit
      -- CP-element group 948: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/SplitProtocol/Sample/ra
      -- 
    ra_9398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 948_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3833_inst_ack_0, ack => zeropad3D_CP_676_elements(948)); -- 
    -- CP-element group 949:  transition  input  bypass 
    -- CP-element group 949: predecessors 
    -- CP-element group 949: 	561 
    -- CP-element group 949: successors 
    -- CP-element group 949: 	950 
    -- CP-element group 949:  members (2) 
      -- CP-element group 949: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/SplitProtocol/Update/$exit
      -- CP-element group 949: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/SplitProtocol/Update/ca
      -- 
    ca_9403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 949_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3833_inst_ack_1, ack => zeropad3D_CP_676_elements(949)); -- 
    -- CP-element group 950:  join  transition  output  bypass 
    -- CP-element group 950: predecessors 
    -- CP-element group 950: 	948 
    -- CP-element group 950: 	949 
    -- CP-element group 950: successors 
    -- CP-element group 950: 	951 
    -- CP-element group 950:  members (5) 
      -- CP-element group 950: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/$exit
      -- CP-element group 950: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/$exit
      -- CP-element group 950: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/$exit
      -- CP-element group 950: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3833/SplitProtocol/$exit
      -- CP-element group 950: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/phi_stmt_3828/phi_stmt_3828_req
      -- 
    phi_stmt_3828_req_9404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3828_req_9404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(950), ack => phi_stmt_3828_req_1); -- 
    zeropad3D_cp_element_group_950: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_950"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(948) & zeropad3D_CP_676_elements(949);
      gj_zeropad3D_cp_element_group_950 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(950), clk => clk, reset => reset); --
    end block;
    -- CP-element group 951:  join  transition  bypass 
    -- CP-element group 951: predecessors 
    -- CP-element group 951: 	944 
    -- CP-element group 951: 	947 
    -- CP-element group 951: 	950 
    -- CP-element group 951: successors 
    -- CP-element group 951: 	952 
    -- CP-element group 951:  members (1) 
      -- CP-element group 951: 	 branch_block_stmt_223/ifx_xthen1744_ifx_xend1784_PhiReq/$exit
      -- 
    zeropad3D_cp_element_group_951: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_951"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(944) & zeropad3D_CP_676_elements(947) & zeropad3D_CP_676_elements(950);
      gj_zeropad3D_cp_element_group_951 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(951), clk => clk, reset => reset); --
    end block;
    -- CP-element group 952:  merge  fork  transition  place  bypass 
    -- CP-element group 952: predecessors 
    -- CP-element group 952: 	941 
    -- CP-element group 952: 	951 
    -- CP-element group 952: successors 
    -- CP-element group 952: 	953 
    -- CP-element group 952: 	954 
    -- CP-element group 952: 	955 
    -- CP-element group 952:  members (2) 
      -- CP-element group 952: 	 branch_block_stmt_223/merge_stmt_3814_PhiReqMerge
      -- CP-element group 952: 	 branch_block_stmt_223/merge_stmt_3814_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(952) <= OrReduce(zeropad3D_CP_676_elements(941) & zeropad3D_CP_676_elements(951));
    -- CP-element group 953:  transition  input  bypass 
    -- CP-element group 953: predecessors 
    -- CP-element group 953: 	952 
    -- CP-element group 953: successors 
    -- CP-element group 953: 	956 
    -- CP-element group 953:  members (1) 
      -- CP-element group 953: 	 branch_block_stmt_223/merge_stmt_3814_PhiAck/phi_stmt_3815_ack
      -- 
    phi_stmt_3815_ack_9409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 953_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3815_ack_0, ack => zeropad3D_CP_676_elements(953)); -- 
    -- CP-element group 954:  transition  input  bypass 
    -- CP-element group 954: predecessors 
    -- CP-element group 954: 	952 
    -- CP-element group 954: successors 
    -- CP-element group 954: 	956 
    -- CP-element group 954:  members (1) 
      -- CP-element group 954: 	 branch_block_stmt_223/merge_stmt_3814_PhiAck/phi_stmt_3822_ack
      -- 
    phi_stmt_3822_ack_9410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 954_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3822_ack_0, ack => zeropad3D_CP_676_elements(954)); -- 
    -- CP-element group 955:  transition  input  bypass 
    -- CP-element group 955: predecessors 
    -- CP-element group 955: 	952 
    -- CP-element group 955: successors 
    -- CP-element group 955: 	956 
    -- CP-element group 955:  members (1) 
      -- CP-element group 955: 	 branch_block_stmt_223/merge_stmt_3814_PhiAck/phi_stmt_3828_ack
      -- 
    phi_stmt_3828_ack_9411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 955_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3828_ack_0, ack => zeropad3D_CP_676_elements(955)); -- 
    -- CP-element group 956:  join  transition  bypass 
    -- CP-element group 956: predecessors 
    -- CP-element group 956: 	953 
    -- CP-element group 956: 	954 
    -- CP-element group 956: 	955 
    -- CP-element group 956: successors 
    -- CP-element group 956: 	8 
    -- CP-element group 956:  members (1) 
      -- CP-element group 956: 	 branch_block_stmt_223/merge_stmt_3814_PhiAck/$exit
      -- 
    zeropad3D_cp_element_group_956: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_956"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(953) & zeropad3D_CP_676_elements(954) & zeropad3D_CP_676_elements(955);
      gj_zeropad3D_cp_element_group_956 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(956), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1165_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1248_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1273_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1579_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1662_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1687_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1977_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2060_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2085_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2393_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2476_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2501_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2791_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2874_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2899_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3195_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3278_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3303_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3605_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3688_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3713_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_555_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_617_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_755_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_839_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_864_wire : std_logic_vector(31 downto 0);
    signal LOAD_pad_1000_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_1000_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_1408_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_1408_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_1813_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_1813_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_2216_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_2216_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_2627_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_2627_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_3030_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_3030_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_3441_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_3441_word_address_0 : std_logic_vector(0 downto 0);
    signal LOAD_pad_512_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_pad_512_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom1023_2404_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1023_2404_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1066_2487_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1066_2487_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1071_2512_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1071_2512_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1246_2802_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1246_2802_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1289_2885_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1289_2885_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1294_2910_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1294_2910_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1464_3206_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1464_3206_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1507_3289_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1507_3289_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1512_3314_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1512_3314_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom157_767_resized : std_logic_vector(13 downto 0);
    signal R_idxprom157_767_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1684_3616_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1684_3616_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1727_3699_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1727_3699_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom1732_3724_resized : std_logic_vector(13 downto 0);
    signal R_idxprom1732_3724_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom197_850_resized : std_logic_vector(13 downto 0);
    signal R_idxprom197_850_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom202_875_resized : std_logic_vector(13 downto 0);
    signal R_idxprom202_875_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom367_1176_resized : std_logic_vector(13 downto 0);
    signal R_idxprom367_1176_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom410_1259_resized : std_logic_vector(13 downto 0);
    signal R_idxprom410_1259_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom415_1284_resized : std_logic_vector(13 downto 0);
    signal R_idxprom415_1284_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom584_1590_resized : std_logic_vector(13 downto 0);
    signal R_idxprom584_1590_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom627_1673_resized : std_logic_vector(13 downto 0);
    signal R_idxprom627_1673_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom632_1698_resized : std_logic_vector(13 downto 0);
    signal R_idxprom632_1698_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom805_1988_resized : std_logic_vector(13 downto 0);
    signal R_idxprom805_1988_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom848_2071_resized : std_logic_vector(13 downto 0);
    signal R_idxprom848_2071_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom853_2096_resized : std_logic_vector(13 downto 0);
    signal R_idxprom853_2096_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_349_resized : std_logic_vector(13 downto 0);
    signal R_indvar_349_scaled : std_logic_vector(13 downto 0);
    signal STORE_pad_242_data_0 : std_logic_vector(7 downto 0);
    signal STORE_pad_242_word_address_0 : std_logic_vector(0 downto 0);
    signal add1001_2259 : std_logic_vector(31 downto 0);
    signal add1014_2381 : std_logic_vector(31 downto 0);
    signal add1020_2386 : std_logic_vector(31 downto 0);
    signal add1038_2444 : std_logic_vector(31 downto 0);
    signal add1047_2449 : std_logic_vector(31 downto 0);
    signal add1057_2464 : std_logic_vector(31 downto 0);
    signal add1063_2469 : std_logic_vector(31 downto 0);
    signal add1078_2532 : std_logic_vector(31 downto 0);
    signal add1086_2552 : std_logic_vector(15 downto 0);
    signal add1099_2232 : std_logic_vector(31 downto 0);
    signal add1116_2249 : std_logic_vector(31 downto 0);
    signal add119_594 : std_logic_vector(31 downto 0);
    signal add1207_2653 : std_logic_vector(31 downto 0);
    signal add1224_2658 : std_logic_vector(31 downto 0);
    signal add1237_2779 : std_logic_vector(31 downto 0);
    signal add1243_2784 : std_logic_vector(31 downto 0);
    signal add1261_2842 : std_logic_vector(31 downto 0);
    signal add1270_2847 : std_logic_vector(31 downto 0);
    signal add1280_2862 : std_logic_vector(31 downto 0);
    signal add1286_2867 : std_logic_vector(31 downto 0);
    signal add1301_2930 : std_logic_vector(31 downto 0);
    signal add1309_2950 : std_logic_vector(15 downto 0);
    signal add1321_2643 : std_logic_vector(31 downto 0);
    signal add1338_2648 : std_logic_vector(31 downto 0);
    signal add137_599 : std_logic_vector(31 downto 0);
    signal add1424_3056 : std_logic_vector(31 downto 0);
    signal add1442_3061 : std_logic_vector(31 downto 0);
    signal add1455_3183 : std_logic_vector(31 downto 0);
    signal add1461_3188 : std_logic_vector(31 downto 0);
    signal add1479_3246 : std_logic_vector(31 downto 0);
    signal add1488_3251 : std_logic_vector(31 downto 0);
    signal add148_743 : std_logic_vector(31 downto 0);
    signal add1498_3266 : std_logic_vector(31 downto 0);
    signal add1504_3271 : std_logic_vector(31 downto 0);
    signal add1519_3334 : std_logic_vector(31 downto 0);
    signal add1527_3354 : std_logic_vector(15 downto 0);
    signal add1540_3046 : std_logic_vector(31 downto 0);
    signal add154_748 : std_logic_vector(31 downto 0);
    signal add1555_3051 : std_logic_vector(31 downto 0);
    signal add1645_3467 : std_logic_vector(31 downto 0);
    signal add1662_3472 : std_logic_vector(31 downto 0);
    signal add1675_3593 : std_logic_vector(31 downto 0);
    signal add1681_3598 : std_logic_vector(31 downto 0);
    signal add1699_3656 : std_logic_vector(31 downto 0);
    signal add169_807 : std_logic_vector(31 downto 0);
    signal add1708_3661 : std_logic_vector(31 downto 0);
    signal add1718_3676 : std_logic_vector(31 downto 0);
    signal add1724_3681 : std_logic_vector(31 downto 0);
    signal add1739_3744 : std_logic_vector(31 downto 0);
    signal add1747_3764 : std_logic_vector(15 downto 0);
    signal add1759_3457 : std_logic_vector(31 downto 0);
    signal add1774_3462 : std_logic_vector(31 downto 0);
    signal add178_812 : std_logic_vector(31 downto 0);
    signal add188_827 : std_logic_vector(31 downto 0);
    signal add194_832 : std_logic_vector(31 downto 0);
    signal add207_895 : std_logic_vector(31 downto 0);
    signal add215_915 : std_logic_vector(15 downto 0);
    signal add228_574 : std_logic_vector(31 downto 0);
    signal add244_589 : std_logic_vector(31 downto 0);
    signal add31_395 : std_logic_vector(63 downto 0);
    signal add328_1026 : std_logic_vector(31 downto 0);
    signal add345_1031 : std_logic_vector(31 downto 0);
    signal add358_1153 : std_logic_vector(31 downto 0);
    signal add364_1158 : std_logic_vector(31 downto 0);
    signal add37_413 : std_logic_vector(63 downto 0);
    signal add382_1216 : std_logic_vector(31 downto 0);
    signal add391_1221 : std_logic_vector(31 downto 0);
    signal add401_1236 : std_logic_vector(31 downto 0);
    signal add407_1241 : std_logic_vector(31 downto 0);
    signal add422_1304 : std_logic_vector(31 downto 0);
    signal add430_1324 : std_logic_vector(15 downto 0);
    signal add43_431 : std_logic_vector(63 downto 0);
    signal add442_1016 : std_logic_vector(31 downto 0);
    signal add458_1021 : std_logic_vector(31 downto 0);
    signal add49_449 : std_logic_vector(63 downto 0);
    signal add544_1440 : std_logic_vector(31 downto 0);
    signal add55_467 : std_logic_vector(63 downto 0);
    signal add562_1445 : std_logic_vector(31 downto 0);
    signal add575_1567 : std_logic_vector(31 downto 0);
    signal add581_1572 : std_logic_vector(31 downto 0);
    signal add599_1630 : std_logic_vector(31 downto 0);
    signal add608_1635 : std_logic_vector(31 downto 0);
    signal add618_1650 : std_logic_vector(31 downto 0);
    signal add61_485 : std_logic_vector(63 downto 0);
    signal add624_1655 : std_logic_vector(31 downto 0);
    signal add639_1718 : std_logic_vector(31 downto 0);
    signal add647_1738 : std_logic_vector(15 downto 0);
    signal add660_1424 : std_logic_vector(31 downto 0);
    signal add676_1435 : std_logic_vector(31 downto 0);
    signal add766_1839 : std_logic_vector(31 downto 0);
    signal add783_1844 : std_logic_vector(31 downto 0);
    signal add796_1965 : std_logic_vector(31 downto 0);
    signal add802_1970 : std_logic_vector(31 downto 0);
    signal add820_2028 : std_logic_vector(31 downto 0);
    signal add829_2033 : std_logic_vector(31 downto 0);
    signal add839_2048 : std_logic_vector(31 downto 0);
    signal add845_2053 : std_logic_vector(31 downto 0);
    signal add860_2116 : std_logic_vector(31 downto 0);
    signal add868_2136 : std_logic_vector(15 downto 0);
    signal add880_1829 : std_logic_vector(31 downto 0);
    signal add896_1834 : std_logic_vector(31 downto 0);
    signal add983_2254 : std_logic_vector(31 downto 0);
    signal add_377 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1177_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1177_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1177_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1177_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1177_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1177_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1260_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1285_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1285_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1285_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1285_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1285_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1285_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1591_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1591_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1591_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1591_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1591_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1591_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1674_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1674_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1674_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1674_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1674_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1674_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1699_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1699_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1699_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1699_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1699_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1699_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1989_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1989_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1989_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1989_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1989_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1989_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2072_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2097_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2405_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2405_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2405_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2405_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2405_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2405_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2488_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2488_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2488_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2488_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2488_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2488_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2513_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2513_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2513_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2513_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2513_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2513_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2803_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2803_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2803_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2803_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2803_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2803_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2886_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2886_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2886_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2886_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2886_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2886_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2911_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2911_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2911_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2911_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2911_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2911_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3207_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3207_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3207_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3207_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3207_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3207_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3290_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3290_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3290_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3290_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3290_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3290_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3315_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3315_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3315_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3315_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3315_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3315_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_350_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3617_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3617_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3617_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3617_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3617_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3617_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3700_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3700_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3700_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3700_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3700_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3700_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_768_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_768_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_768_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_768_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_768_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_768_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_851_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_851_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_851_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_851_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_851_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_851_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_root_address : std_logic_vector(13 downto 0);
    signal arrayidx1024_2407 : std_logic_vector(31 downto 0);
    signal arrayidx1067_2490 : std_logic_vector(31 downto 0);
    signal arrayidx1072_2515 : std_logic_vector(31 downto 0);
    signal arrayidx1247_2805 : std_logic_vector(31 downto 0);
    signal arrayidx1290_2888 : std_logic_vector(31 downto 0);
    signal arrayidx1295_2913 : std_logic_vector(31 downto 0);
    signal arrayidx1465_3209 : std_logic_vector(31 downto 0);
    signal arrayidx1508_3292 : std_logic_vector(31 downto 0);
    signal arrayidx1513_3317 : std_logic_vector(31 downto 0);
    signal arrayidx158_770 : std_logic_vector(31 downto 0);
    signal arrayidx1685_3619 : std_logic_vector(31 downto 0);
    signal arrayidx1728_3702 : std_logic_vector(31 downto 0);
    signal arrayidx1733_3727 : std_logic_vector(31 downto 0);
    signal arrayidx198_853 : std_logic_vector(31 downto 0);
    signal arrayidx203_878 : std_logic_vector(31 downto 0);
    signal arrayidx368_1179 : std_logic_vector(31 downto 0);
    signal arrayidx411_1262 : std_logic_vector(31 downto 0);
    signal arrayidx416_1287 : std_logic_vector(31 downto 0);
    signal arrayidx585_1593 : std_logic_vector(31 downto 0);
    signal arrayidx628_1676 : std_logic_vector(31 downto 0);
    signal arrayidx633_1701 : std_logic_vector(31 downto 0);
    signal arrayidx806_1991 : std_logic_vector(31 downto 0);
    signal arrayidx849_2074 : std_logic_vector(31 downto 0);
    signal arrayidx854_2099 : std_logic_vector(31 downto 0);
    signal arrayidx_352 : std_logic_vector(31 downto 0);
    signal call1_229 : std_logic_vector(7 downto 0);
    signal call20_355 : std_logic_vector(7 downto 0);
    signal call23_368 : std_logic_vector(7 downto 0);
    signal call28_386 : std_logic_vector(7 downto 0);
    signal call2_232 : std_logic_vector(7 downto 0);
    signal call34_404 : std_logic_vector(7 downto 0);
    signal call3_235 : std_logic_vector(7 downto 0);
    signal call40_422 : std_logic_vector(7 downto 0);
    signal call46_440 : std_logic_vector(7 downto 0);
    signal call4_238 : std_logic_vector(7 downto 0);
    signal call52_458 : std_logic_vector(7 downto 0);
    signal call58_476 : std_logic_vector(7 downto 0);
    signal call5_241 : std_logic_vector(7 downto 0);
    signal call6_247 : std_logic_vector(7 downto 0);
    signal call7_250 : std_logic_vector(7 downto 0);
    signal call8_253 : std_logic_vector(7 downto 0);
    signal call_226 : std_logic_vector(7 downto 0);
    signal cmp1002_2344 : std_logic_vector(0 downto 0);
    signal cmp1081_2539 : std_logic_vector(0 downto 0);
    signal cmp1100_2570 : std_logic_vector(0 downto 0);
    signal cmp1117_2596 : std_logic_vector(0 downto 0);
    signal cmp111_656 : std_logic_vector(0 downto 0);
    signal cmp111x_xnot_662 : std_logic_vector(0 downto 0);
    signal cmp1196_2692 : std_logic_vector(0 downto 0);
    signal cmp1196x_xnot_2698 : std_logic_vector(0 downto 0);
    signal cmp1208_2705 : std_logic_vector(0 downto 0);
    signal cmp120_669 : std_logic_vector(0 downto 0);
    signal cmp1215_2729 : std_logic_vector(0 downto 0);
    signal cmp1215x_xnot_2735 : std_logic_vector(0 downto 0);
    signal cmp1225_2742 : std_logic_vector(0 downto 0);
    signal cmp127_693 : std_logic_vector(0 downto 0);
    signal cmp127x_xnot_699 : std_logic_vector(0 downto 0);
    signal cmp1304_2937 : std_logic_vector(0 downto 0);
    signal cmp1322_2968 : std_logic_vector(0 downto 0);
    signal cmp1339_2993 : std_logic_vector(0 downto 0);
    signal cmp138_706 : std_logic_vector(0 downto 0);
    signal cmp1415_3096 : std_logic_vector(0 downto 0);
    signal cmp1415x_xnot_3102 : std_logic_vector(0 downto 0);
    signal cmp1425_3109 : std_logic_vector(0 downto 0);
    signal cmp1432_3133 : std_logic_vector(0 downto 0);
    signal cmp1432x_xnot_3139 : std_logic_vector(0 downto 0);
    signal cmp1443_3146 : std_logic_vector(0 downto 0);
    signal cmp1522_3341 : std_logic_vector(0 downto 0);
    signal cmp1541_3372 : std_logic_vector(0 downto 0);
    signal cmp1556_3398 : std_logic_vector(0 downto 0);
    signal cmp1636_3506 : std_logic_vector(0 downto 0);
    signal cmp1636x_xnot_3512 : std_logic_vector(0 downto 0);
    signal cmp1646_3519 : std_logic_vector(0 downto 0);
    signal cmp1653_3543 : std_logic_vector(0 downto 0);
    signal cmp1653x_xnot_3549 : std_logic_vector(0 downto 0);
    signal cmp1663_3556 : std_logic_vector(0 downto 0);
    signal cmp1742_3751 : std_logic_vector(0 downto 0);
    signal cmp1760_3782 : std_logic_vector(0 downto 0);
    signal cmp1775_3807 : std_logic_vector(0 downto 0);
    signal cmp1840_287 : std_logic_vector(0 downto 0);
    signal cmp210_902 : std_logic_vector(0 downto 0);
    signal cmp229_933 : std_logic_vector(0 downto 0);
    signal cmp245_959 : std_logic_vector(0 downto 0);
    signal cmp318_1066 : std_logic_vector(0 downto 0);
    signal cmp318x_xnot_1072 : std_logic_vector(0 downto 0);
    signal cmp329_1079 : std_logic_vector(0 downto 0);
    signal cmp336_1103 : std_logic_vector(0 downto 0);
    signal cmp336x_xnot_1109 : std_logic_vector(0 downto 0);
    signal cmp346_1116 : std_logic_vector(0 downto 0);
    signal cmp425_1311 : std_logic_vector(0 downto 0);
    signal cmp443_1342 : std_logic_vector(0 downto 0);
    signal cmp459_1367 : std_logic_vector(0 downto 0);
    signal cmp534_1480 : std_logic_vector(0 downto 0);
    signal cmp534x_xnot_1486 : std_logic_vector(0 downto 0);
    signal cmp545_1493 : std_logic_vector(0 downto 0);
    signal cmp552_1517 : std_logic_vector(0 downto 0);
    signal cmp552x_xnot_1523 : std_logic_vector(0 downto 0);
    signal cmp563_1530 : std_logic_vector(0 downto 0);
    signal cmp642_1725 : std_logic_vector(0 downto 0);
    signal cmp661_1756 : std_logic_vector(0 downto 0);
    signal cmp677_1782 : std_logic_vector(0 downto 0);
    signal cmp756_1878 : std_logic_vector(0 downto 0);
    signal cmp756x_xnot_1884 : std_logic_vector(0 downto 0);
    signal cmp767_1891 : std_logic_vector(0 downto 0);
    signal cmp774_1915 : std_logic_vector(0 downto 0);
    signal cmp774x_xnot_1921 : std_logic_vector(0 downto 0);
    signal cmp784_1928 : std_logic_vector(0 downto 0);
    signal cmp863_2123 : std_logic_vector(0 downto 0);
    signal cmp881_2154 : std_logic_vector(0 downto 0);
    signal cmp897_2179 : std_logic_vector(0 downto 0);
    signal cmp972_2294 : std_logic_vector(0 downto 0);
    signal cmp972x_xnot_2300 : std_logic_vector(0 downto 0);
    signal cmp984_2307 : std_logic_vector(0 downto 0);
    signal cmp991_2331 : std_logic_vector(0 downto 0);
    signal cmp991x_xnot_2337 : std_logic_vector(0 downto 0);
    signal conv1008_2361 : std_logic_vector(31 downto 0);
    signal conv1012_2366 : std_logic_vector(31 downto 0);
    signal conv101_529 : std_logic_vector(31 downto 0);
    signal conv1029_2419 : std_logic_vector(31 downto 0);
    signal conv1077_2526 : std_logic_vector(31 downto 0);
    signal conv108_649 : std_logic_vector(31 downto 0);
    signal conv1092_2565 : std_logic_vector(31 downto 0);
    signal conv10_261 : std_logic_vector(63 downto 0);
    signal conv1108_2591 : std_logic_vector(31 downto 0);
    signal conv110_538 : std_logic_vector(31 downto 0);
    signal conv1193_2685 : std_logic_vector(31 downto 0);
    signal conv1195_2632 : std_logic_vector(31 downto 0);
    signal conv1212_2722 : std_logic_vector(31 downto 0);
    signal conv1231_2759 : std_logic_vector(31 downto 0);
    signal conv1235_2764 : std_logic_vector(31 downto 0);
    signal conv124_686 : std_logic_vector(31 downto 0);
    signal conv1252_2817 : std_logic_vector(31 downto 0);
    signal conv12_265 : std_logic_vector(63 downto 0);
    signal conv1300_2924 : std_logic_vector(31 downto 0);
    signal conv1315_2963 : std_logic_vector(31 downto 0);
    signal conv1330_2988 : std_logic_vector(31 downto 0);
    signal conv1412_3089 : std_logic_vector(31 downto 0);
    signal conv1414_3035 : std_logic_vector(31 downto 0);
    signal conv1429_3126 : std_logic_vector(31 downto 0);
    signal conv142_723 : std_logic_vector(31 downto 0);
    signal conv1449_3163 : std_logic_vector(31 downto 0);
    signal conv144_542 : std_logic_vector(31 downto 0);
    signal conv1453_3168 : std_logic_vector(31 downto 0);
    signal conv146_728 : std_logic_vector(31 downto 0);
    signal conv1470_3221 : std_logic_vector(31 downto 0);
    signal conv150_557 : std_logic_vector(31 downto 0);
    signal conv1518_3328 : std_logic_vector(31 downto 0);
    signal conv1533_3367 : std_logic_vector(31 downto 0);
    signal conv1549_3393 : std_logic_vector(31 downto 0);
    signal conv161_782 : std_logic_vector(31 downto 0);
    signal conv1633_3499 : std_logic_vector(31 downto 0);
    signal conv1635_3446 : std_logic_vector(31 downto 0);
    signal conv1650_3536 : std_logic_vector(31 downto 0);
    signal conv1669_3573 : std_logic_vector(31 downto 0);
    signal conv1673_3578 : std_logic_vector(31 downto 0);
    signal conv1690_3631 : std_logic_vector(31 downto 0);
    signal conv171_619 : std_logic_vector(31 downto 0);
    signal conv1738_3738 : std_logic_vector(31 downto 0);
    signal conv1753_3777 : std_logic_vector(31 downto 0);
    signal conv1768_3802 : std_logic_vector(31 downto 0);
    signal conv1788_3841 : std_logic_vector(31 downto 0);
    signal conv1790_3845 : std_logic_vector(31 downto 0);
    signal conv206_889 : std_logic_vector(31 downto 0);
    signal conv21_359 : std_logic_vector(63 downto 0);
    signal conv221_928 : std_logic_vector(31 downto 0);
    signal conv237_954 : std_logic_vector(31 downto 0);
    signal conv239_578 : std_logic_vector(31 downto 0);
    signal conv259_992 : std_logic_vector(15 downto 0);
    signal conv25_372 : std_logic_vector(63 downto 0);
    signal conv30_390 : std_logic_vector(63 downto 0);
    signal conv315_1059 : std_logic_vector(31 downto 0);
    signal conv317_1005 : std_logic_vector(31 downto 0);
    signal conv333_1096 : std_logic_vector(31 downto 0);
    signal conv352_1133 : std_logic_vector(31 downto 0);
    signal conv356_1138 : std_logic_vector(31 downto 0);
    signal conv36_408 : std_logic_vector(63 downto 0);
    signal conv373_1191 : std_logic_vector(31 downto 0);
    signal conv421_1298 : std_logic_vector(31 downto 0);
    signal conv42_426 : std_logic_vector(63 downto 0);
    signal conv436_1337 : std_logic_vector(31 downto 0);
    signal conv451_1362 : std_logic_vector(31 downto 0);
    signal conv477_1400 : std_logic_vector(15 downto 0);
    signal conv48_444 : std_logic_vector(63 downto 0);
    signal conv531_1473 : std_logic_vector(31 downto 0);
    signal conv533_1413 : std_logic_vector(31 downto 0);
    signal conv549_1510 : std_logic_vector(31 downto 0);
    signal conv54_462 : std_logic_vector(63 downto 0);
    signal conv569_1547 : std_logic_vector(31 downto 0);
    signal conv573_1552 : std_logic_vector(31 downto 0);
    signal conv590_1605 : std_logic_vector(31 downto 0);
    signal conv60_480 : std_logic_vector(63 downto 0);
    signal conv638_1712 : std_logic_vector(31 downto 0);
    signal conv653_1751 : std_logic_vector(31 downto 0);
    signal conv669_1777 : std_logic_vector(31 downto 0);
    signal conv753_1871 : std_logic_vector(31 downto 0);
    signal conv755_1818 : std_logic_vector(31 downto 0);
    signal conv771_1908 : std_logic_vector(31 downto 0);
    signal conv790_1945 : std_logic_vector(31 downto 0);
    signal conv794_1950 : std_logic_vector(31 downto 0);
    signal conv811_2003 : std_logic_vector(31 downto 0);
    signal conv859_2110 : std_logic_vector(31 downto 0);
    signal conv874_2149 : std_logic_vector(31 downto 0);
    signal conv889_2174 : std_logic_vector(31 downto 0);
    signal conv92_517 : std_logic_vector(31 downto 0);
    signal conv94_521 : std_logic_vector(31 downto 0);
    signal conv969_2287 : std_logic_vector(31 downto 0);
    signal conv971_2221 : std_logic_vector(31 downto 0);
    signal conv988_2324 : std_logic_vector(31 downto 0);
    signal conv99_525 : std_logic_vector(31 downto 0);
    signal conv_257 : std_logic_vector(63 downto 0);
    signal div1112_2244 : std_logic_vector(31 downto 0);
    signal div1580_3439 : std_logic_vector(15 downto 0);
    signal div224_563 : std_logic_vector(31 downto 0);
    signal div240_584 : std_logic_vector(31 downto 0);
    signal div260_998 : std_logic_vector(15 downto 0);
    signal div478_1406 : std_logic_vector(15 downto 0);
    signal div672_1430 : std_logic_vector(31 downto 0);
    signal div916_2214 : std_logic_vector(15 downto 0);
    signal exitcond8_500 : std_logic_vector(0 downto 0);
    signal i1137x_x1x_xph_3008 : std_logic_vector(15 downto 0);
    signal i1137x_x2_2668 : std_logic_vector(15 downto 0);
    signal i1355x_x1x_xph_3413 : std_logic_vector(15 downto 0);
    signal i1355x_x2_3071 : std_logic_vector(15 downto 0);
    signal i1576x_x1x_xph_3822 : std_logic_vector(15 downto 0);
    signal i1576x_x2_3482 : std_logic_vector(15 downto 0);
    signal i263x_x1x_xph_1381 : std_logic_vector(15 downto 0);
    signal i263x_x2_1040 : std_logic_vector(15 downto 0);
    signal i475x_x1x_xph_1797 : std_logic_vector(15 downto 0);
    signal i475x_x2_1455 : std_logic_vector(15 downto 0);
    signal i68x_x1x_xph_973 : std_logic_vector(15 downto 0);
    signal i68x_x2_630 : std_logic_vector(15 downto 0);
    signal i697x_x1x_xph_2194 : std_logic_vector(15 downto 0);
    signal i697x_x2_1854 : std_logic_vector(15 downto 0);
    signal i913x_x1x_xph_2611 : std_logic_vector(15 downto 0);
    signal i913x_x2_2269 : std_logic_vector(15 downto 0);
    signal idxprom1023_2400 : std_logic_vector(63 downto 0);
    signal idxprom1066_2483 : std_logic_vector(63 downto 0);
    signal idxprom1071_2508 : std_logic_vector(63 downto 0);
    signal idxprom1246_2798 : std_logic_vector(63 downto 0);
    signal idxprom1289_2881 : std_logic_vector(63 downto 0);
    signal idxprom1294_2906 : std_logic_vector(63 downto 0);
    signal idxprom1464_3202 : std_logic_vector(63 downto 0);
    signal idxprom1507_3285 : std_logic_vector(63 downto 0);
    signal idxprom1512_3310 : std_logic_vector(63 downto 0);
    signal idxprom157_763 : std_logic_vector(63 downto 0);
    signal idxprom1684_3612 : std_logic_vector(63 downto 0);
    signal idxprom1727_3695 : std_logic_vector(63 downto 0);
    signal idxprom1732_3720 : std_logic_vector(63 downto 0);
    signal idxprom197_846 : std_logic_vector(63 downto 0);
    signal idxprom202_871 : std_logic_vector(63 downto 0);
    signal idxprom367_1172 : std_logic_vector(63 downto 0);
    signal idxprom410_1255 : std_logic_vector(63 downto 0);
    signal idxprom415_1280 : std_logic_vector(63 downto 0);
    signal idxprom584_1586 : std_logic_vector(63 downto 0);
    signal idxprom627_1669 : std_logic_vector(63 downto 0);
    signal idxprom632_1694 : std_logic_vector(63 downto 0);
    signal idxprom805_1984 : std_logic_vector(63 downto 0);
    signal idxprom848_2067 : std_logic_vector(63 downto 0);
    signal idxprom853_2092 : std_logic_vector(63 downto 0);
    signal inc1090_2560 : std_logic_vector(15 downto 0);
    signal inc1105_2574 : std_logic_vector(15 downto 0);
    signal inc1105x_xi913x_x2_2579 : std_logic_vector(15 downto 0);
    signal inc1313_2958 : std_logic_vector(15 downto 0);
    signal inc1327_2972 : std_logic_vector(15 downto 0);
    signal inc1327x_xi1137x_x2_2977 : std_logic_vector(15 downto 0);
    signal inc1531_3362 : std_logic_vector(15 downto 0);
    signal inc1546_3376 : std_logic_vector(15 downto 0);
    signal inc1546x_xi1355x_x2_3381 : std_logic_vector(15 downto 0);
    signal inc1751_3772 : std_logic_vector(15 downto 0);
    signal inc1765_3786 : std_logic_vector(15 downto 0);
    signal inc1765x_xi1576x_x2_3791 : std_logic_vector(15 downto 0);
    signal inc219_923 : std_logic_vector(15 downto 0);
    signal inc234_937 : std_logic_vector(15 downto 0);
    signal inc234x_xi68x_x2_942 : std_logic_vector(15 downto 0);
    signal inc434_1332 : std_logic_vector(15 downto 0);
    signal inc448_1346 : std_logic_vector(15 downto 0);
    signal inc448x_xi263x_x2_1351 : std_logic_vector(15 downto 0);
    signal inc651_1746 : std_logic_vector(15 downto 0);
    signal inc666_1760 : std_logic_vector(15 downto 0);
    signal inc666x_xi475x_x2_1765 : std_logic_vector(15 downto 0);
    signal inc872_2144 : std_logic_vector(15 downto 0);
    signal inc886_2158 : std_logic_vector(15 downto 0);
    signal inc886x_xi697x_x2_2163 : std_logic_vector(15 downto 0);
    signal indvar_338 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_495 : std_logic_vector(63 downto 0);
    signal j1187x_x0x_xph_3014 : std_logic_vector(15 downto 0);
    signal j1187x_x1_2674 : std_logic_vector(15 downto 0);
    signal j1187x_x2_2983 : std_logic_vector(15 downto 0);
    signal j1406x_x0x_xph_3419 : std_logic_vector(15 downto 0);
    signal j1406x_x1_3077 : std_logic_vector(15 downto 0);
    signal j1406x_x2_3388 : std_logic_vector(15 downto 0);
    signal j1627x_x0x_xph_3828 : std_logic_vector(15 downto 0);
    signal j1627x_x1_3488 : std_logic_vector(15 downto 0);
    signal j1627x_x2_3797 : std_logic_vector(15 downto 0);
    signal j309x_x0x_xph_1375 : std_logic_vector(15 downto 0);
    signal j309x_x1_1034 : std_logic_vector(15 downto 0);
    signal j309x_x2_1357 : std_logic_vector(15 downto 0);
    signal j525x_x0x_xph_1803 : std_logic_vector(15 downto 0);
    signal j525x_x1_1461 : std_logic_vector(15 downto 0);
    signal j525x_x2_1772 : std_logic_vector(15 downto 0);
    signal j747x_x0x_xph_2200 : std_logic_vector(15 downto 0);
    signal j747x_x1_1860 : std_logic_vector(15 downto 0);
    signal j747x_x2_2169 : std_logic_vector(15 downto 0);
    signal j963x_x0x_xph_2617 : std_logic_vector(15 downto 0);
    signal j963x_x1_2275 : std_logic_vector(15 downto 0);
    signal j963x_x2_2586 : std_logic_vector(15 downto 0);
    signal jx_x0x_xph_967 : std_logic_vector(15 downto 0);
    signal jx_x1_622 : std_logic_vector(15 downto 0);
    signal jx_x2_949 : std_logic_vector(15 downto 0);
    signal k1129x_x0x_xph_3001 : std_logic_vector(15 downto 0);
    signal k1129x_x1_2661 : std_logic_vector(15 downto 0);
    signal k1351x_x0x_xph_3406 : std_logic_vector(15 downto 0);
    signal k1351x_x1_3064 : std_logic_vector(15 downto 0);
    signal k1568x_x0x_xph_3815 : std_logic_vector(15 downto 0);
    signal k1568x_x1_3475 : std_logic_vector(15 downto 0);
    signal k255x_x0x_xph_1387 : std_logic_vector(15 downto 0);
    signal k255x_x1_1047 : std_logic_vector(15 downto 0);
    signal k471x_x0x_xph_1790 : std_logic_vector(15 downto 0);
    signal k471x_x1_1448 : std_logic_vector(15 downto 0);
    signal k689x_x0x_xph_2187 : std_logic_vector(15 downto 0);
    signal k689x_x1_1847 : std_logic_vector(15 downto 0);
    signal k909x_x0x_xph_2604 : std_logic_vector(15 downto 0);
    signal k909x_x1_2262 : std_logic_vector(15 downto 0);
    signal kx_x0x_xph_979 : std_logic_vector(15 downto 0);
    signal kx_x1_637 : std_logic_vector(15 downto 0);
    signal mul1013_2371 : std_logic_vector(31 downto 0);
    signal mul1019_2376 : std_logic_vector(31 downto 0);
    signal mul102_534 : std_logic_vector(31 downto 0);
    signal mul1037_2429 : std_logic_vector(31 downto 0);
    signal mul1046_2439 : std_logic_vector(31 downto 0);
    signal mul1056_2454 : std_logic_vector(31 downto 0);
    signal mul1062_2459 : std_logic_vector(31 downto 0);
    signal mul1111_2238 : std_logic_vector(31 downto 0);
    signal mul1236_2769 : std_logic_vector(31 downto 0);
    signal mul1242_2774 : std_logic_vector(31 downto 0);
    signal mul1260_2827 : std_logic_vector(31 downto 0);
    signal mul1269_2837 : std_logic_vector(31 downto 0);
    signal mul1279_2852 : std_logic_vector(31 downto 0);
    signal mul1285_2857 : std_logic_vector(31 downto 0);
    signal mul1359_3028 : std_logic_vector(15 downto 0);
    signal mul13_275 : std_logic_vector(63 downto 0);
    signal mul1454_3173 : std_logic_vector(31 downto 0);
    signal mul1460_3178 : std_logic_vector(31 downto 0);
    signal mul1478_3231 : std_logic_vector(31 downto 0);
    signal mul147_733 : std_logic_vector(31 downto 0);
    signal mul1487_3241 : std_logic_vector(31 downto 0);
    signal mul1497_3256 : std_logic_vector(31 downto 0);
    signal mul1503_3261 : std_logic_vector(31 downto 0);
    signal mul153_738 : std_logic_vector(31 downto 0);
    signal mul1579_3433 : std_logic_vector(15 downto 0);
    signal mul1674_3583 : std_logic_vector(31 downto 0);
    signal mul1680_3588 : std_logic_vector(31 downto 0);
    signal mul168_792 : std_logic_vector(31 downto 0);
    signal mul1698_3641 : std_logic_vector(31 downto 0);
    signal mul1707_3651 : std_logic_vector(31 downto 0);
    signal mul1717_3666 : std_logic_vector(31 downto 0);
    signal mul1723_3671 : std_logic_vector(31 downto 0);
    signal mul177_802 : std_logic_vector(31 downto 0);
    signal mul1791_3850 : std_logic_vector(31 downto 0);
    signal mul1794_3855 : std_logic_vector(31 downto 0);
    signal mul187_817 : std_logic_vector(31 downto 0);
    signal mul193_822 : std_logic_vector(31 downto 0);
    signal mul357_1143 : std_logic_vector(31 downto 0);
    signal mul363_1148 : std_logic_vector(31 downto 0);
    signal mul381_1201 : std_logic_vector(31 downto 0);
    signal mul390_1211 : std_logic_vector(31 downto 0);
    signal mul400_1226 : std_logic_vector(31 downto 0);
    signal mul406_1231 : std_logic_vector(31 downto 0);
    signal mul574_1557 : std_logic_vector(31 downto 0);
    signal mul580_1562 : std_logic_vector(31 downto 0);
    signal mul598_1615 : std_logic_vector(31 downto 0);
    signal mul607_1625 : std_logic_vector(31 downto 0);
    signal mul617_1640 : std_logic_vector(31 downto 0);
    signal mul623_1645 : std_logic_vector(31 downto 0);
    signal mul795_1955 : std_logic_vector(31 downto 0);
    signal mul801_1960 : std_logic_vector(31 downto 0);
    signal mul819_2013 : std_logic_vector(31 downto 0);
    signal mul828_2023 : std_logic_vector(31 downto 0);
    signal mul838_2038 : std_logic_vector(31 downto 0);
    signal mul844_2043 : std_logic_vector(31 downto 0);
    signal mul95_605 : std_logic_vector(31 downto 0);
    signal mul_270 : std_logic_vector(63 downto 0);
    signal orx_xcond1849_711 : std_logic_vector(0 downto 0);
    signal orx_xcond1850_1084 : std_logic_vector(0 downto 0);
    signal orx_xcond1851_1121 : std_logic_vector(0 downto 0);
    signal orx_xcond1852_1498 : std_logic_vector(0 downto 0);
    signal orx_xcond1853_1535 : std_logic_vector(0 downto 0);
    signal orx_xcond1854_1896 : std_logic_vector(0 downto 0);
    signal orx_xcond1855_1933 : std_logic_vector(0 downto 0);
    signal orx_xcond1856_2312 : std_logic_vector(0 downto 0);
    signal orx_xcond1857_2349 : std_logic_vector(0 downto 0);
    signal orx_xcond1858_2710 : std_logic_vector(0 downto 0);
    signal orx_xcond1859_2747 : std_logic_vector(0 downto 0);
    signal orx_xcond1860_3114 : std_logic_vector(0 downto 0);
    signal orx_xcond1861_3151 : std_logic_vector(0 downto 0);
    signal orx_xcond1862_3524 : std_logic_vector(0 downto 0);
    signal orx_xcond1863_3561 : std_logic_vector(0 downto 0);
    signal orx_xcond_674 : std_logic_vector(0 downto 0);
    signal ptr_deref_1181_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1181_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1181_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1181_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1181_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1181_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1265_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1265_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1265_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1265_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1265_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1289_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1289_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1289_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1289_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1289_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1289_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1595_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1595_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1595_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1595_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1595_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1595_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1679_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1679_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1679_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1679_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1679_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1703_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1703_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1703_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1703_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1703_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1703_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1993_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1993_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1993_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1993_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1993_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1993_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2077_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2077_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2077_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2077_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2077_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2101_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2101_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2101_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2101_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2101_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2101_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2409_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2409_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2409_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2409_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2409_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2409_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2493_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2493_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2493_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2493_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2493_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2517_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2517_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2517_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2517_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2517_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2517_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2807_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2807_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2807_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2807_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2807_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2807_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2891_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2891_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2891_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2891_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2891_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2915_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2915_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2915_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2915_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2915_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2915_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3211_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3211_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3211_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3211_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3211_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3211_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3295_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3295_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3295_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3295_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3295_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3319_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3319_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3319_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3319_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3319_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3319_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3621_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3621_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3621_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3621_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3621_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3621_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3705_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3705_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3705_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3705_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3705_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3729_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3729_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3729_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3729_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3729_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3729_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_487_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_487_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_487_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_487_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_487_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_487_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_772_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_772_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_772_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_772_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_772_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_772_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_856_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_856_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_856_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_856_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_856_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_880_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_880_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_880_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_880_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_880_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_880_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext1848_548 : std_logic_vector(31 downto 0);
    signal sext_610 : std_logic_vector(31 downto 0);
    signal shl1098_2227 : std_logic_vector(31 downto 0);
    signal shl1320_2638 : std_logic_vector(31 downto 0);
    signal shl1539_3041 : std_logic_vector(31 downto 0);
    signal shl1758_3452 : std_logic_vector(31 downto 0);
    signal shl227_569 : std_logic_vector(31 downto 0);
    signal shl27_383 : std_logic_vector(63 downto 0);
    signal shl33_401 : std_logic_vector(63 downto 0);
    signal shl39_419 : std_logic_vector(63 downto 0);
    signal shl441_1011 : std_logic_vector(31 downto 0);
    signal shl45_437 : std_logic_vector(63 downto 0);
    signal shl51_455 : std_logic_vector(63 downto 0);
    signal shl57_473 : std_logic_vector(63 downto 0);
    signal shl659_1419 : std_logic_vector(31 downto 0);
    signal shl879_1824 : std_logic_vector(31 downto 0);
    signal shl_365 : std_logic_vector(63 downto 0);
    signal shr1022_2395 : std_logic_vector(31 downto 0);
    signal shr1065_2478 : std_logic_vector(31 downto 0);
    signal shr1070_2503 : std_logic_vector(31 downto 0);
    signal shr1245_2793 : std_logic_vector(31 downto 0);
    signal shr1288_2876 : std_logic_vector(31 downto 0);
    signal shr1293_2901 : std_logic_vector(31 downto 0);
    signal shr1463_3197 : std_logic_vector(31 downto 0);
    signal shr1506_3280 : std_logic_vector(31 downto 0);
    signal shr1511_3305 : std_logic_vector(31 downto 0);
    signal shr156_757 : std_logic_vector(31 downto 0);
    signal shr1683_3607 : std_logic_vector(31 downto 0);
    signal shr1726_3690 : std_logic_vector(31 downto 0);
    signal shr1731_3715 : std_logic_vector(31 downto 0);
    signal shr1839x_xmask_281 : std_logic_vector(63 downto 0);
    signal shr196_841 : std_logic_vector(31 downto 0);
    signal shr201_866 : std_logic_vector(31 downto 0);
    signal shr366_1167 : std_logic_vector(31 downto 0);
    signal shr409_1250 : std_logic_vector(31 downto 0);
    signal shr414_1275 : std_logic_vector(31 downto 0);
    signal shr583_1581 : std_logic_vector(31 downto 0);
    signal shr626_1664 : std_logic_vector(31 downto 0);
    signal shr631_1689 : std_logic_vector(31 downto 0);
    signal shr804_1979 : std_logic_vector(31 downto 0);
    signal shr847_2062 : std_logic_vector(31 downto 0);
    signal shr852_2087 : std_logic_vector(31 downto 0);
    signal sub1036_2424 : std_logic_vector(31 downto 0);
    signal sub1045_2434 : std_logic_vector(31 downto 0);
    signal sub1259_2822 : std_logic_vector(31 downto 0);
    signal sub1268_2832 : std_logic_vector(31 downto 0);
    signal sub1477_3226 : std_logic_vector(31 downto 0);
    signal sub1486_3236 : std_logic_vector(31 downto 0);
    signal sub1697_3636 : std_logic_vector(31 downto 0);
    signal sub1706_3646 : std_logic_vector(31 downto 0);
    signal sub176_797 : std_logic_vector(31 downto 0);
    signal sub380_1196 : std_logic_vector(31 downto 0);
    signal sub389_1206 : std_logic_vector(31 downto 0);
    signal sub597_1610 : std_logic_vector(31 downto 0);
    signal sub606_1620 : std_logic_vector(31 downto 0);
    signal sub818_2008 : std_logic_vector(31 downto 0);
    signal sub827_2018 : std_logic_vector(31 downto 0);
    signal sub_787 : std_logic_vector(31 downto 0);
    signal tmp1068_2494 : std_logic_vector(63 downto 0);
    signal tmp1144_2628 : std_logic_vector(7 downto 0);
    signal tmp1291_2892 : std_logic_vector(63 downto 0);
    signal tmp1363_3031 : std_logic_vector(7 downto 0);
    signal tmp1509_3296 : std_logic_vector(63 downto 0);
    signal tmp1584_3442 : std_logic_vector(7 downto 0);
    signal tmp1729_3706 : std_logic_vector(63 downto 0);
    signal tmp199_857 : std_logic_vector(63 downto 0);
    signal tmp1_302 : std_logic_vector(63 downto 0);
    signal tmp266_1001 : std_logic_vector(7 downto 0);
    signal tmp2_307 : std_logic_vector(63 downto 0);
    signal tmp3_311 : std_logic_vector(63 downto 0);
    signal tmp412_1266 : std_logic_vector(63 downto 0);
    signal tmp482_1409 : std_logic_vector(7 downto 0);
    signal tmp4_316 : std_logic_vector(63 downto 0);
    signal tmp5_322 : std_logic_vector(63 downto 0);
    signal tmp629_1680 : std_logic_vector(63 downto 0);
    signal tmp6_328 : std_logic_vector(0 downto 0);
    signal tmp704_1814 : std_logic_vector(7 downto 0);
    signal tmp70_513 : std_logic_vector(7 downto 0);
    signal tmp850_2078 : std_logic_vector(63 downto 0);
    signal tmp920_2217 : std_logic_vector(7 downto 0);
    signal tmp_298 : std_logic_vector(63 downto 0);
    signal type_cast_1009_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1037_wire : std_logic_vector(15 downto 0);
    signal type_cast_1039_wire : std_logic_vector(15 downto 0);
    signal type_cast_1044_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1046_wire : std_logic_vector(15 downto 0);
    signal type_cast_1051_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1053_wire : std_logic_vector(15 downto 0);
    signal type_cast_1057_wire : std_logic_vector(31 downto 0);
    signal type_cast_1062_wire : std_logic_vector(31 downto 0);
    signal type_cast_1064_wire : std_logic_vector(31 downto 0);
    signal type_cast_1070_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1075_wire : std_logic_vector(31 downto 0);
    signal type_cast_1077_wire : std_logic_vector(31 downto 0);
    signal type_cast_1094_wire : std_logic_vector(31 downto 0);
    signal type_cast_1099_wire : std_logic_vector(31 downto 0);
    signal type_cast_1101_wire : std_logic_vector(31 downto 0);
    signal type_cast_1107_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1112_wire : std_logic_vector(31 downto 0);
    signal type_cast_1114_wire : std_logic_vector(31 downto 0);
    signal type_cast_1131_wire : std_logic_vector(31 downto 0);
    signal type_cast_1136_wire : std_logic_vector(31 downto 0);
    signal type_cast_1161_wire : std_logic_vector(31 downto 0);
    signal type_cast_1164_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1170_wire : std_logic_vector(63 downto 0);
    signal type_cast_1183_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1189_wire : std_logic_vector(31 downto 0);
    signal type_cast_1244_wire : std_logic_vector(31 downto 0);
    signal type_cast_1247_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1253_wire : std_logic_vector(63 downto 0);
    signal type_cast_1269_wire : std_logic_vector(31 downto 0);
    signal type_cast_1272_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1278_wire : std_logic_vector(63 downto 0);
    signal type_cast_1296_wire : std_logic_vector(31 downto 0);
    signal type_cast_1302_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1307_wire : std_logic_vector(31 downto 0);
    signal type_cast_1309_wire : std_logic_vector(31 downto 0);
    signal type_cast_1322_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1330_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1335_wire : std_logic_vector(31 downto 0);
    signal type_cast_1360_wire : std_logic_vector(31 downto 0);
    signal type_cast_1378_wire : std_logic_vector(15 downto 0);
    signal type_cast_1380_wire : std_logic_vector(15 downto 0);
    signal type_cast_1384_wire : std_logic_vector(15 downto 0);
    signal type_cast_1386_wire : std_logic_vector(15 downto 0);
    signal type_cast_1390_wire : std_logic_vector(15 downto 0);
    signal type_cast_1393_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1404_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1417_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1428_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1452_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1454_wire : std_logic_vector(15 downto 0);
    signal type_cast_1458_wire : std_logic_vector(15 downto 0);
    signal type_cast_1460_wire : std_logic_vector(15 downto 0);
    signal type_cast_1465_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1467_wire : std_logic_vector(15 downto 0);
    signal type_cast_1471_wire : std_logic_vector(31 downto 0);
    signal type_cast_1476_wire : std_logic_vector(31 downto 0);
    signal type_cast_1478_wire : std_logic_vector(31 downto 0);
    signal type_cast_1484_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1489_wire : std_logic_vector(31 downto 0);
    signal type_cast_1491_wire : std_logic_vector(31 downto 0);
    signal type_cast_1508_wire : std_logic_vector(31 downto 0);
    signal type_cast_1513_wire : std_logic_vector(31 downto 0);
    signal type_cast_1515_wire : std_logic_vector(31 downto 0);
    signal type_cast_1521_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1526_wire : std_logic_vector(31 downto 0);
    signal type_cast_1528_wire : std_logic_vector(31 downto 0);
    signal type_cast_1545_wire : std_logic_vector(31 downto 0);
    signal type_cast_1550_wire : std_logic_vector(31 downto 0);
    signal type_cast_1575_wire : std_logic_vector(31 downto 0);
    signal type_cast_1578_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1584_wire : std_logic_vector(63 downto 0);
    signal type_cast_1597_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1603_wire : std_logic_vector(31 downto 0);
    signal type_cast_1658_wire : std_logic_vector(31 downto 0);
    signal type_cast_1661_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1667_wire : std_logic_vector(63 downto 0);
    signal type_cast_1683_wire : std_logic_vector(31 downto 0);
    signal type_cast_1686_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1692_wire : std_logic_vector(63 downto 0);
    signal type_cast_1710_wire : std_logic_vector(31 downto 0);
    signal type_cast_1716_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1721_wire : std_logic_vector(31 downto 0);
    signal type_cast_1723_wire : std_logic_vector(31 downto 0);
    signal type_cast_1736_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1744_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1749_wire : std_logic_vector(31 downto 0);
    signal type_cast_1769_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1775_wire : std_logic_vector(31 downto 0);
    signal type_cast_1793_wire : std_logic_vector(15 downto 0);
    signal type_cast_1796_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1800_wire : std_logic_vector(15 downto 0);
    signal type_cast_1802_wire : std_logic_vector(15 downto 0);
    signal type_cast_1806_wire : std_logic_vector(15 downto 0);
    signal type_cast_1808_wire : std_logic_vector(15 downto 0);
    signal type_cast_1822_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1850_wire : std_logic_vector(15 downto 0);
    signal type_cast_1853_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1857_wire : std_logic_vector(15 downto 0);
    signal type_cast_1859_wire : std_logic_vector(15 downto 0);
    signal type_cast_1863_wire : std_logic_vector(15 downto 0);
    signal type_cast_1865_wire : std_logic_vector(15 downto 0);
    signal type_cast_1869_wire : std_logic_vector(31 downto 0);
    signal type_cast_1874_wire : std_logic_vector(31 downto 0);
    signal type_cast_1876_wire : std_logic_vector(31 downto 0);
    signal type_cast_1882_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1887_wire : std_logic_vector(31 downto 0);
    signal type_cast_1889_wire : std_logic_vector(31 downto 0);
    signal type_cast_1906_wire : std_logic_vector(31 downto 0);
    signal type_cast_1911_wire : std_logic_vector(31 downto 0);
    signal type_cast_1913_wire : std_logic_vector(31 downto 0);
    signal type_cast_1919_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1924_wire : std_logic_vector(31 downto 0);
    signal type_cast_1926_wire : std_logic_vector(31 downto 0);
    signal type_cast_1943_wire : std_logic_vector(31 downto 0);
    signal type_cast_1948_wire : std_logic_vector(31 downto 0);
    signal type_cast_1973_wire : std_logic_vector(31 downto 0);
    signal type_cast_1976_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1982_wire : std_logic_vector(63 downto 0);
    signal type_cast_1995_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2001_wire : std_logic_vector(31 downto 0);
    signal type_cast_2056_wire : std_logic_vector(31 downto 0);
    signal type_cast_2059_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2065_wire : std_logic_vector(63 downto 0);
    signal type_cast_2081_wire : std_logic_vector(31 downto 0);
    signal type_cast_2084_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2090_wire : std_logic_vector(63 downto 0);
    signal type_cast_2108_wire : std_logic_vector(31 downto 0);
    signal type_cast_2114_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2119_wire : std_logic_vector(31 downto 0);
    signal type_cast_2121_wire : std_logic_vector(31 downto 0);
    signal type_cast_2134_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2142_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2147_wire : std_logic_vector(31 downto 0);
    signal type_cast_2172_wire : std_logic_vector(31 downto 0);
    signal type_cast_2191_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2193_wire : std_logic_vector(15 downto 0);
    signal type_cast_2197_wire : std_logic_vector(15 downto 0);
    signal type_cast_2199_wire : std_logic_vector(15 downto 0);
    signal type_cast_2203_wire : std_logic_vector(15 downto 0);
    signal type_cast_2205_wire : std_logic_vector(15 downto 0);
    signal type_cast_2212_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2225_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2236_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2242_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2266_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2268_wire : std_logic_vector(15 downto 0);
    signal type_cast_2272_wire : std_logic_vector(15 downto 0);
    signal type_cast_2274_wire : std_logic_vector(15 downto 0);
    signal type_cast_2279_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2281_wire : std_logic_vector(15 downto 0);
    signal type_cast_2285_wire : std_logic_vector(31 downto 0);
    signal type_cast_2290_wire : std_logic_vector(31 downto 0);
    signal type_cast_2292_wire : std_logic_vector(31 downto 0);
    signal type_cast_2298_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2303_wire : std_logic_vector(31 downto 0);
    signal type_cast_2305_wire : std_logic_vector(31 downto 0);
    signal type_cast_2322_wire : std_logic_vector(31 downto 0);
    signal type_cast_2327_wire : std_logic_vector(31 downto 0);
    signal type_cast_2329_wire : std_logic_vector(31 downto 0);
    signal type_cast_2335_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2340_wire : std_logic_vector(31 downto 0);
    signal type_cast_2342_wire : std_logic_vector(31 downto 0);
    signal type_cast_2359_wire : std_logic_vector(31 downto 0);
    signal type_cast_2364_wire : std_logic_vector(31 downto 0);
    signal type_cast_2389_wire : std_logic_vector(31 downto 0);
    signal type_cast_2392_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2398_wire : std_logic_vector(63 downto 0);
    signal type_cast_2411_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2417_wire : std_logic_vector(31 downto 0);
    signal type_cast_2472_wire : std_logic_vector(31 downto 0);
    signal type_cast_2475_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2481_wire : std_logic_vector(63 downto 0);
    signal type_cast_2497_wire : std_logic_vector(31 downto 0);
    signal type_cast_2500_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2506_wire : std_logic_vector(63 downto 0);
    signal type_cast_2524_wire : std_logic_vector(31 downto 0);
    signal type_cast_2530_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2535_wire : std_logic_vector(31 downto 0);
    signal type_cast_2537_wire : std_logic_vector(31 downto 0);
    signal type_cast_2550_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2558_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2563_wire : std_logic_vector(31 downto 0);
    signal type_cast_2583_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2589_wire : std_logic_vector(31 downto 0);
    signal type_cast_2607_wire : std_logic_vector(15 downto 0);
    signal type_cast_2610_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2614_wire : std_logic_vector(15 downto 0);
    signal type_cast_2616_wire : std_logic_vector(15 downto 0);
    signal type_cast_2620_wire : std_logic_vector(15 downto 0);
    signal type_cast_2622_wire : std_logic_vector(15 downto 0);
    signal type_cast_2636_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2665_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2667_wire : std_logic_vector(15 downto 0);
    signal type_cast_2671_wire : std_logic_vector(15 downto 0);
    signal type_cast_2673_wire : std_logic_vector(15 downto 0);
    signal type_cast_2677_wire : std_logic_vector(15 downto 0);
    signal type_cast_2679_wire : std_logic_vector(15 downto 0);
    signal type_cast_2683_wire : std_logic_vector(31 downto 0);
    signal type_cast_2688_wire : std_logic_vector(31 downto 0);
    signal type_cast_2690_wire : std_logic_vector(31 downto 0);
    signal type_cast_2696_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2701_wire : std_logic_vector(31 downto 0);
    signal type_cast_2703_wire : std_logic_vector(31 downto 0);
    signal type_cast_2720_wire : std_logic_vector(31 downto 0);
    signal type_cast_2725_wire : std_logic_vector(31 downto 0);
    signal type_cast_2727_wire : std_logic_vector(31 downto 0);
    signal type_cast_2733_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2738_wire : std_logic_vector(31 downto 0);
    signal type_cast_2740_wire : std_logic_vector(31 downto 0);
    signal type_cast_2757_wire : std_logic_vector(31 downto 0);
    signal type_cast_2762_wire : std_logic_vector(31 downto 0);
    signal type_cast_2787_wire : std_logic_vector(31 downto 0);
    signal type_cast_2790_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2796_wire : std_logic_vector(63 downto 0);
    signal type_cast_279_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2809_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2815_wire : std_logic_vector(31 downto 0);
    signal type_cast_285_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2870_wire : std_logic_vector(31 downto 0);
    signal type_cast_2873_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2879_wire : std_logic_vector(63 downto 0);
    signal type_cast_2895_wire : std_logic_vector(31 downto 0);
    signal type_cast_2898_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2904_wire : std_logic_vector(63 downto 0);
    signal type_cast_2922_wire : std_logic_vector(31 downto 0);
    signal type_cast_2928_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2933_wire : std_logic_vector(31 downto 0);
    signal type_cast_2935_wire : std_logic_vector(31 downto 0);
    signal type_cast_2948_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2956_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2961_wire : std_logic_vector(31 downto 0);
    signal type_cast_2986_wire : std_logic_vector(31 downto 0);
    signal type_cast_3004_wire : std_logic_vector(15 downto 0);
    signal type_cast_3007_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3011_wire : std_logic_vector(15 downto 0);
    signal type_cast_3013_wire : std_logic_vector(15 downto 0);
    signal type_cast_3017_wire : std_logic_vector(15 downto 0);
    signal type_cast_3019_wire : std_logic_vector(15 downto 0);
    signal type_cast_3026_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3039_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3068_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3070_wire : std_logic_vector(15 downto 0);
    signal type_cast_3074_wire : std_logic_vector(15 downto 0);
    signal type_cast_3076_wire : std_logic_vector(15 downto 0);
    signal type_cast_3080_wire : std_logic_vector(15 downto 0);
    signal type_cast_3083_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3087_wire : std_logic_vector(31 downto 0);
    signal type_cast_3092_wire : std_logic_vector(31 downto 0);
    signal type_cast_3094_wire : std_logic_vector(31 downto 0);
    signal type_cast_3100_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3105_wire : std_logic_vector(31 downto 0);
    signal type_cast_3107_wire : std_logic_vector(31 downto 0);
    signal type_cast_3124_wire : std_logic_vector(31 downto 0);
    signal type_cast_3129_wire : std_logic_vector(31 downto 0);
    signal type_cast_3131_wire : std_logic_vector(31 downto 0);
    signal type_cast_3137_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3142_wire : std_logic_vector(31 downto 0);
    signal type_cast_3144_wire : std_logic_vector(31 downto 0);
    signal type_cast_3161_wire : std_logic_vector(31 downto 0);
    signal type_cast_3166_wire : std_logic_vector(31 downto 0);
    signal type_cast_3191_wire : std_logic_vector(31 downto 0);
    signal type_cast_3194_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3200_wire : std_logic_vector(63 downto 0);
    signal type_cast_320_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3213_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3219_wire : std_logic_vector(31 downto 0);
    signal type_cast_326_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3274_wire : std_logic_vector(31 downto 0);
    signal type_cast_3277_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3283_wire : std_logic_vector(63 downto 0);
    signal type_cast_3299_wire : std_logic_vector(31 downto 0);
    signal type_cast_3302_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3308_wire : std_logic_vector(63 downto 0);
    signal type_cast_3326_wire : std_logic_vector(31 downto 0);
    signal type_cast_3332_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3337_wire : std_logic_vector(31 downto 0);
    signal type_cast_3339_wire : std_logic_vector(31 downto 0);
    signal type_cast_333_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3352_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3360_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3365_wire : std_logic_vector(31 downto 0);
    signal type_cast_3385_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3391_wire : std_logic_vector(31 downto 0);
    signal type_cast_3410_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3412_wire : std_logic_vector(15 downto 0);
    signal type_cast_3416_wire : std_logic_vector(15 downto 0);
    signal type_cast_3418_wire : std_logic_vector(15 downto 0);
    signal type_cast_3422_wire : std_logic_vector(15 downto 0);
    signal type_cast_3424_wire : std_logic_vector(15 downto 0);
    signal type_cast_342_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3431_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3437_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_344_wire : std_logic_vector(63 downto 0);
    signal type_cast_3450_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3479_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3481_wire : std_logic_vector(15 downto 0);
    signal type_cast_3485_wire : std_logic_vector(15 downto 0);
    signal type_cast_3487_wire : std_logic_vector(15 downto 0);
    signal type_cast_3491_wire : std_logic_vector(15 downto 0);
    signal type_cast_3493_wire : std_logic_vector(15 downto 0);
    signal type_cast_3497_wire : std_logic_vector(31 downto 0);
    signal type_cast_3502_wire : std_logic_vector(31 downto 0);
    signal type_cast_3504_wire : std_logic_vector(31 downto 0);
    signal type_cast_3510_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3515_wire : std_logic_vector(31 downto 0);
    signal type_cast_3517_wire : std_logic_vector(31 downto 0);
    signal type_cast_3534_wire : std_logic_vector(31 downto 0);
    signal type_cast_3539_wire : std_logic_vector(31 downto 0);
    signal type_cast_3541_wire : std_logic_vector(31 downto 0);
    signal type_cast_3547_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3552_wire : std_logic_vector(31 downto 0);
    signal type_cast_3554_wire : std_logic_vector(31 downto 0);
    signal type_cast_3571_wire : std_logic_vector(31 downto 0);
    signal type_cast_3576_wire : std_logic_vector(31 downto 0);
    signal type_cast_3601_wire : std_logic_vector(31 downto 0);
    signal type_cast_3604_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3610_wire : std_logic_vector(63 downto 0);
    signal type_cast_3623_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3629_wire : std_logic_vector(31 downto 0);
    signal type_cast_363_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3684_wire : std_logic_vector(31 downto 0);
    signal type_cast_3687_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3693_wire : std_logic_vector(63 downto 0);
    signal type_cast_3709_wire : std_logic_vector(31 downto 0);
    signal type_cast_3712_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3718_wire : std_logic_vector(63 downto 0);
    signal type_cast_3736_wire : std_logic_vector(31 downto 0);
    signal type_cast_3742_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3747_wire : std_logic_vector(31 downto 0);
    signal type_cast_3749_wire : std_logic_vector(31 downto 0);
    signal type_cast_3762_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3770_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3775_wire : std_logic_vector(31 downto 0);
    signal type_cast_3800_wire : std_logic_vector(31 downto 0);
    signal type_cast_3819_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_381_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3821_wire : std_logic_vector(15 downto 0);
    signal type_cast_3825_wire : std_logic_vector(15 downto 0);
    signal type_cast_3827_wire : std_logic_vector(15 downto 0);
    signal type_cast_3831_wire : std_logic_vector(15 downto 0);
    signal type_cast_3833_wire : std_logic_vector(15 downto 0);
    signal type_cast_399_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_417_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_435_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_453_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_471_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_493_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_546_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_551_wire : std_logic_vector(31 downto 0);
    signal type_cast_554_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_561_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_567_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_582_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_603_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_613_wire : std_logic_vector(31 downto 0);
    signal type_cast_616_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_627_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_629_wire : std_logic_vector(15 downto 0);
    signal type_cast_634_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_636_wire : std_logic_vector(15 downto 0);
    signal type_cast_641_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_643_wire : std_logic_vector(15 downto 0);
    signal type_cast_647_wire : std_logic_vector(31 downto 0);
    signal type_cast_652_wire : std_logic_vector(31 downto 0);
    signal type_cast_654_wire : std_logic_vector(31 downto 0);
    signal type_cast_660_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_665_wire : std_logic_vector(31 downto 0);
    signal type_cast_667_wire : std_logic_vector(31 downto 0);
    signal type_cast_684_wire : std_logic_vector(31 downto 0);
    signal type_cast_689_wire : std_logic_vector(31 downto 0);
    signal type_cast_691_wire : std_logic_vector(31 downto 0);
    signal type_cast_697_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_702_wire : std_logic_vector(31 downto 0);
    signal type_cast_704_wire : std_logic_vector(31 downto 0);
    signal type_cast_721_wire : std_logic_vector(31 downto 0);
    signal type_cast_726_wire : std_logic_vector(31 downto 0);
    signal type_cast_751_wire : std_logic_vector(31 downto 0);
    signal type_cast_754_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_761_wire : std_logic_vector(63 downto 0);
    signal type_cast_774_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_780_wire : std_logic_vector(31 downto 0);
    signal type_cast_835_wire : std_logic_vector(31 downto 0);
    signal type_cast_838_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_844_wire : std_logic_vector(63 downto 0);
    signal type_cast_860_wire : std_logic_vector(31 downto 0);
    signal type_cast_863_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_869_wire : std_logic_vector(63 downto 0);
    signal type_cast_887_wire : std_logic_vector(31 downto 0);
    signal type_cast_893_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_898_wire : std_logic_vector(31 downto 0);
    signal type_cast_900_wire : std_logic_vector(31 downto 0);
    signal type_cast_913_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_921_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_926_wire : std_logic_vector(31 downto 0);
    signal type_cast_946_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_952_wire : std_logic_vector(31 downto 0);
    signal type_cast_970_wire : std_logic_vector(15 downto 0);
    signal type_cast_972_wire : std_logic_vector(15 downto 0);
    signal type_cast_976_wire : std_logic_vector(15 downto 0);
    signal type_cast_978_wire : std_logic_vector(15 downto 0);
    signal type_cast_982_wire : std_logic_vector(15 downto 0);
    signal type_cast_985_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_996_wire_constant : std_logic_vector(15 downto 0);
    signal umax7_335 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    LOAD_pad_1000_word_address_0 <= "0";
    LOAD_pad_1408_word_address_0 <= "0";
    LOAD_pad_1813_word_address_0 <= "0";
    LOAD_pad_2216_word_address_0 <= "0";
    LOAD_pad_2627_word_address_0 <= "0";
    LOAD_pad_3030_word_address_0 <= "0";
    LOAD_pad_3441_word_address_0 <= "0";
    LOAD_pad_512_word_address_0 <= "0";
    STORE_pad_242_word_address_0 <= "0";
    array_obj_ref_1177_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1177_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1177_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1177_resized_base_address <= "00000000000000";
    array_obj_ref_1260_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1260_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1260_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1260_resized_base_address <= "00000000000000";
    array_obj_ref_1285_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1285_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1285_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1285_resized_base_address <= "00000000000000";
    array_obj_ref_1591_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1591_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1591_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1591_resized_base_address <= "00000000000000";
    array_obj_ref_1674_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1674_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1674_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1674_resized_base_address <= "00000000000000";
    array_obj_ref_1699_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1699_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1699_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1699_resized_base_address <= "00000000000000";
    array_obj_ref_1989_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1989_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1989_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1989_resized_base_address <= "00000000000000";
    array_obj_ref_2072_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2072_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2072_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2072_resized_base_address <= "00000000000000";
    array_obj_ref_2097_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2097_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2097_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2097_resized_base_address <= "00000000000000";
    array_obj_ref_2405_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2405_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2405_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2405_resized_base_address <= "00000000000000";
    array_obj_ref_2488_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2488_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2488_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2488_resized_base_address <= "00000000000000";
    array_obj_ref_2513_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2513_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2513_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2513_resized_base_address <= "00000000000000";
    array_obj_ref_2803_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2803_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2803_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2803_resized_base_address <= "00000000000000";
    array_obj_ref_2886_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2886_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2886_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2886_resized_base_address <= "00000000000000";
    array_obj_ref_2911_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2911_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2911_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2911_resized_base_address <= "00000000000000";
    array_obj_ref_3207_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3207_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3207_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3207_resized_base_address <= "00000000000000";
    array_obj_ref_3290_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3290_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3290_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3290_resized_base_address <= "00000000000000";
    array_obj_ref_3315_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3315_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3315_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3315_resized_base_address <= "00000000000000";
    array_obj_ref_350_constant_part_of_offset <= "00000000000000";
    array_obj_ref_350_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_350_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_350_resized_base_address <= "00000000000000";
    array_obj_ref_3617_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3617_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3617_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3617_resized_base_address <= "00000000000000";
    array_obj_ref_3700_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3700_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3700_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3700_resized_base_address <= "00000000000000";
    array_obj_ref_3725_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3725_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3725_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3725_resized_base_address <= "00000000000000";
    array_obj_ref_768_constant_part_of_offset <= "00000000000000";
    array_obj_ref_768_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_768_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_768_resized_base_address <= "00000000000000";
    array_obj_ref_851_constant_part_of_offset <= "00000000000000";
    array_obj_ref_851_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_851_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_851_resized_base_address <= "00000000000000";
    array_obj_ref_876_constant_part_of_offset <= "00000000000000";
    array_obj_ref_876_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_876_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_876_resized_base_address <= "00000000000000";
    ptr_deref_1181_word_offset_0 <= "00000000000000";
    ptr_deref_1265_word_offset_0 <= "00000000000000";
    ptr_deref_1289_word_offset_0 <= "00000000000000";
    ptr_deref_1595_word_offset_0 <= "00000000000000";
    ptr_deref_1679_word_offset_0 <= "00000000000000";
    ptr_deref_1703_word_offset_0 <= "00000000000000";
    ptr_deref_1993_word_offset_0 <= "00000000000000";
    ptr_deref_2077_word_offset_0 <= "00000000000000";
    ptr_deref_2101_word_offset_0 <= "00000000000000";
    ptr_deref_2409_word_offset_0 <= "00000000000000";
    ptr_deref_2493_word_offset_0 <= "00000000000000";
    ptr_deref_2517_word_offset_0 <= "00000000000000";
    ptr_deref_2807_word_offset_0 <= "00000000000000";
    ptr_deref_2891_word_offset_0 <= "00000000000000";
    ptr_deref_2915_word_offset_0 <= "00000000000000";
    ptr_deref_3211_word_offset_0 <= "00000000000000";
    ptr_deref_3295_word_offset_0 <= "00000000000000";
    ptr_deref_3319_word_offset_0 <= "00000000000000";
    ptr_deref_3621_word_offset_0 <= "00000000000000";
    ptr_deref_3705_word_offset_0 <= "00000000000000";
    ptr_deref_3729_word_offset_0 <= "00000000000000";
    ptr_deref_487_word_offset_0 <= "00000000000000";
    ptr_deref_772_word_offset_0 <= "00000000000000";
    ptr_deref_856_word_offset_0 <= "00000000000000";
    ptr_deref_880_word_offset_0 <= "00000000000000";
    type_cast_1009_wire_constant <= "00000000000000000000000000000001";
    type_cast_1044_wire_constant <= "0000000000000000";
    type_cast_1051_wire_constant <= "0000000000000000";
    type_cast_1070_wire_constant <= "1";
    type_cast_1107_wire_constant <= "1";
    type_cast_1164_wire_constant <= "00000000000000000000000000000010";
    type_cast_1183_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1247_wire_constant <= "00000000000000000000000000000010";
    type_cast_1272_wire_constant <= "00000000000000000000000000000010";
    type_cast_1302_wire_constant <= "00000000000000000000000000000100";
    type_cast_1322_wire_constant <= "0000000000000100";
    type_cast_1330_wire_constant <= "0000000000000001";
    type_cast_1393_wire_constant <= "0000000000000000";
    type_cast_1404_wire_constant <= "0000000000000010";
    type_cast_1417_wire_constant <= "00000000000000000000000000000001";
    type_cast_1428_wire_constant <= "00000000000000000000000000000001";
    type_cast_1452_wire_constant <= "0000000000000000";
    type_cast_1465_wire_constant <= "0000000000000000";
    type_cast_1484_wire_constant <= "1";
    type_cast_1521_wire_constant <= "1";
    type_cast_1578_wire_constant <= "00000000000000000000000000000010";
    type_cast_1597_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1661_wire_constant <= "00000000000000000000000000000010";
    type_cast_1686_wire_constant <= "00000000000000000000000000000010";
    type_cast_1716_wire_constant <= "00000000000000000000000000000100";
    type_cast_1736_wire_constant <= "0000000000000100";
    type_cast_1744_wire_constant <= "0000000000000001";
    type_cast_1769_wire_constant <= "0000000000000000";
    type_cast_1796_wire_constant <= "0000000000000000";
    type_cast_1822_wire_constant <= "00000000000000000000000000000001";
    type_cast_1853_wire_constant <= "0000000000000000";
    type_cast_1882_wire_constant <= "1";
    type_cast_1919_wire_constant <= "1";
    type_cast_1976_wire_constant <= "00000000000000000000000000000010";
    type_cast_1995_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2059_wire_constant <= "00000000000000000000000000000010";
    type_cast_2084_wire_constant <= "00000000000000000000000000000010";
    type_cast_2114_wire_constant <= "00000000000000000000000000000100";
    type_cast_2134_wire_constant <= "0000000000000100";
    type_cast_2142_wire_constant <= "0000000000000001";
    type_cast_2191_wire_constant <= "0000000000000000";
    type_cast_2212_wire_constant <= "0000000000000001";
    type_cast_2225_wire_constant <= "00000000000000000000000000000001";
    type_cast_2236_wire_constant <= "00000000000000000000000000000011";
    type_cast_2242_wire_constant <= "00000000000000000000000000000010";
    type_cast_2266_wire_constant <= "0000000000000000";
    type_cast_2279_wire_constant <= "0000000000000000";
    type_cast_2298_wire_constant <= "1";
    type_cast_2335_wire_constant <= "1";
    type_cast_2392_wire_constant <= "00000000000000000000000000000010";
    type_cast_2411_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2475_wire_constant <= "00000000000000000000000000000010";
    type_cast_2500_wire_constant <= "00000000000000000000000000000010";
    type_cast_2530_wire_constant <= "00000000000000000000000000000100";
    type_cast_2550_wire_constant <= "0000000000000100";
    type_cast_2558_wire_constant <= "0000000000000001";
    type_cast_2583_wire_constant <= "0000000000000000";
    type_cast_2610_wire_constant <= "0000000000000000";
    type_cast_2636_wire_constant <= "00000000000000000000000000000001";
    type_cast_2665_wire_constant <= "0000000000000000";
    type_cast_2696_wire_constant <= "1";
    type_cast_2733_wire_constant <= "1";
    type_cast_2790_wire_constant <= "00000000000000000000000000000010";
    type_cast_279_wire_constant <= "0000000000000000000000000000000000000000111111111111111111111100";
    type_cast_2809_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_285_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2873_wire_constant <= "00000000000000000000000000000010";
    type_cast_2898_wire_constant <= "00000000000000000000000000000010";
    type_cast_2928_wire_constant <= "00000000000000000000000000000100";
    type_cast_2948_wire_constant <= "0000000000000100";
    type_cast_2956_wire_constant <= "0000000000000001";
    type_cast_3007_wire_constant <= "0000000000000000";
    type_cast_3026_wire_constant <= "0000000000000011";
    type_cast_3039_wire_constant <= "00000000000000000000000000000001";
    type_cast_3068_wire_constant <= "0000000000000000";
    type_cast_3083_wire_constant <= "0000000000000000";
    type_cast_3100_wire_constant <= "1";
    type_cast_3137_wire_constant <= "1";
    type_cast_3194_wire_constant <= "00000000000000000000000000000010";
    type_cast_320_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_3213_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_326_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_3277_wire_constant <= "00000000000000000000000000000010";
    type_cast_3302_wire_constant <= "00000000000000000000000000000010";
    type_cast_3332_wire_constant <= "00000000000000000000000000000100";
    type_cast_333_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_3352_wire_constant <= "0000000000000100";
    type_cast_3360_wire_constant <= "0000000000000001";
    type_cast_3385_wire_constant <= "0000000000000000";
    type_cast_3410_wire_constant <= "0000000000000000";
    type_cast_342_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_3431_wire_constant <= "0000000000000011";
    type_cast_3437_wire_constant <= "0000000000000010";
    type_cast_3450_wire_constant <= "00000000000000000000000000000001";
    type_cast_3479_wire_constant <= "0000000000000000";
    type_cast_3510_wire_constant <= "1";
    type_cast_3547_wire_constant <= "1";
    type_cast_3604_wire_constant <= "00000000000000000000000000000010";
    type_cast_3623_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_363_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_3687_wire_constant <= "00000000000000000000000000000010";
    type_cast_3712_wire_constant <= "00000000000000000000000000000010";
    type_cast_3742_wire_constant <= "00000000000000000000000000000100";
    type_cast_3762_wire_constant <= "0000000000000100";
    type_cast_3770_wire_constant <= "0000000000000001";
    type_cast_3819_wire_constant <= "0000000000000000";
    type_cast_381_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_399_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_417_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_435_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_453_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_471_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_493_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_546_wire_constant <= "00000000000000000000000000010000";
    type_cast_554_wire_constant <= "00000000000000000000000000010000";
    type_cast_561_wire_constant <= "00000000000000000000000000000001";
    type_cast_567_wire_constant <= "00000000000000000000000000000001";
    type_cast_582_wire_constant <= "00000000000000000000000000000010";
    type_cast_603_wire_constant <= "00000000000000000000000000010000";
    type_cast_616_wire_constant <= "00000000000000000000000000010000";
    type_cast_627_wire_constant <= "0000000000000000";
    type_cast_634_wire_constant <= "0000000000000000";
    type_cast_641_wire_constant <= "0000000000000000";
    type_cast_660_wire_constant <= "1";
    type_cast_697_wire_constant <= "1";
    type_cast_754_wire_constant <= "00000000000000000000000000000010";
    type_cast_774_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_838_wire_constant <= "00000000000000000000000000000010";
    type_cast_863_wire_constant <= "00000000000000000000000000000010";
    type_cast_893_wire_constant <= "00000000000000000000000000000100";
    type_cast_913_wire_constant <= "0000000000000100";
    type_cast_921_wire_constant <= "0000000000000001";
    type_cast_946_wire_constant <= "0000000000000000";
    type_cast_985_wire_constant <= "0000000000000000";
    type_cast_996_wire_constant <= "0000000000000001";
    phi_stmt_1034: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1037_wire & type_cast_1039_wire;
      req <= phi_stmt_1034_req_0 & phi_stmt_1034_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1034",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1034_ack_0,
          idata => idata,
          odata => j309x_x1_1034,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1034
    phi_stmt_1040: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1044_wire_constant & type_cast_1046_wire;
      req <= phi_stmt_1040_req_0 & phi_stmt_1040_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1040",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1040_ack_0,
          idata => idata,
          odata => i263x_x2_1040,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1040
    phi_stmt_1047: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1051_wire_constant & type_cast_1053_wire;
      req <= phi_stmt_1047_req_0 & phi_stmt_1047_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1047",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1047_ack_0,
          idata => idata,
          odata => k255x_x1_1047,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1047
    phi_stmt_1375: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1378_wire & type_cast_1380_wire;
      req <= phi_stmt_1375_req_0 & phi_stmt_1375_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1375",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1375_ack_0,
          idata => idata,
          odata => j309x_x0x_xph_1375,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1375
    phi_stmt_1381: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1384_wire & type_cast_1386_wire;
      req <= phi_stmt_1381_req_0 & phi_stmt_1381_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1381",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1381_ack_0,
          idata => idata,
          odata => i263x_x1x_xph_1381,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1381
    phi_stmt_1387: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1390_wire & type_cast_1393_wire_constant;
      req <= phi_stmt_1387_req_0 & phi_stmt_1387_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1387",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1387_ack_0,
          idata => idata,
          odata => k255x_x0x_xph_1387,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1387
    phi_stmt_1448: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1452_wire_constant & type_cast_1454_wire;
      req <= phi_stmt_1448_req_0 & phi_stmt_1448_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1448",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1448_ack_0,
          idata => idata,
          odata => k471x_x1_1448,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1448
    phi_stmt_1455: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1458_wire & type_cast_1460_wire;
      req <= phi_stmt_1455_req_0 & phi_stmt_1455_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1455",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1455_ack_0,
          idata => idata,
          odata => i475x_x2_1455,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1455
    phi_stmt_1461: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1465_wire_constant & type_cast_1467_wire;
      req <= phi_stmt_1461_req_0 & phi_stmt_1461_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1461",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1461_ack_0,
          idata => idata,
          odata => j525x_x1_1461,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1461
    phi_stmt_1790: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1793_wire & type_cast_1796_wire_constant;
      req <= phi_stmt_1790_req_0 & phi_stmt_1790_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1790",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1790_ack_0,
          idata => idata,
          odata => k471x_x0x_xph_1790,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1790
    phi_stmt_1797: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1800_wire & type_cast_1802_wire;
      req <= phi_stmt_1797_req_0 & phi_stmt_1797_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1797",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1797_ack_0,
          idata => idata,
          odata => i475x_x1x_xph_1797,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1797
    phi_stmt_1803: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1806_wire & type_cast_1808_wire;
      req <= phi_stmt_1803_req_0 & phi_stmt_1803_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1803",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1803_ack_0,
          idata => idata,
          odata => j525x_x0x_xph_1803,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1803
    phi_stmt_1847: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1850_wire & type_cast_1853_wire_constant;
      req <= phi_stmt_1847_req_0 & phi_stmt_1847_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1847",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1847_ack_0,
          idata => idata,
          odata => k689x_x1_1847,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1847
    phi_stmt_1854: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1857_wire & type_cast_1859_wire;
      req <= phi_stmt_1854_req_0 & phi_stmt_1854_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1854",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1854_ack_0,
          idata => idata,
          odata => i697x_x2_1854,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1854
    phi_stmt_1860: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1863_wire & type_cast_1865_wire;
      req <= phi_stmt_1860_req_0 & phi_stmt_1860_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1860",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1860_ack_0,
          idata => idata,
          odata => j747x_x1_1860,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1860
    phi_stmt_2187: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2191_wire_constant & type_cast_2193_wire;
      req <= phi_stmt_2187_req_0 & phi_stmt_2187_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2187",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2187_ack_0,
          idata => idata,
          odata => k689x_x0x_xph_2187,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2187
    phi_stmt_2194: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2197_wire & type_cast_2199_wire;
      req <= phi_stmt_2194_req_0 & phi_stmt_2194_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2194",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2194_ack_0,
          idata => idata,
          odata => i697x_x1x_xph_2194,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2194
    phi_stmt_2200: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2203_wire & type_cast_2205_wire;
      req <= phi_stmt_2200_req_0 & phi_stmt_2200_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2200",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2200_ack_0,
          idata => idata,
          odata => j747x_x0x_xph_2200,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2200
    phi_stmt_2262: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2266_wire_constant & type_cast_2268_wire;
      req <= phi_stmt_2262_req_0 & phi_stmt_2262_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2262",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2262_ack_0,
          idata => idata,
          odata => k909x_x1_2262,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2262
    phi_stmt_2269: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2272_wire & type_cast_2274_wire;
      req <= phi_stmt_2269_req_0 & phi_stmt_2269_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2269",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2269_ack_0,
          idata => idata,
          odata => i913x_x2_2269,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2269
    phi_stmt_2275: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2279_wire_constant & type_cast_2281_wire;
      req <= phi_stmt_2275_req_0 & phi_stmt_2275_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2275",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2275_ack_0,
          idata => idata,
          odata => j963x_x1_2275,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2275
    phi_stmt_2604: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2607_wire & type_cast_2610_wire_constant;
      req <= phi_stmt_2604_req_0 & phi_stmt_2604_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2604",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2604_ack_0,
          idata => idata,
          odata => k909x_x0x_xph_2604,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2604
    phi_stmt_2611: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2614_wire & type_cast_2616_wire;
      req <= phi_stmt_2611_req_0 & phi_stmt_2611_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2611",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2611_ack_0,
          idata => idata,
          odata => i913x_x1x_xph_2611,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2611
    phi_stmt_2617: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2620_wire & type_cast_2622_wire;
      req <= phi_stmt_2617_req_0 & phi_stmt_2617_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2617",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2617_ack_0,
          idata => idata,
          odata => j963x_x0x_xph_2617,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2617
    phi_stmt_2661: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2665_wire_constant & type_cast_2667_wire;
      req <= phi_stmt_2661_req_0 & phi_stmt_2661_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2661",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2661_ack_0,
          idata => idata,
          odata => k1129x_x1_2661,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2661
    phi_stmt_2668: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2671_wire & type_cast_2673_wire;
      req <= phi_stmt_2668_req_0 & phi_stmt_2668_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2668",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2668_ack_0,
          idata => idata,
          odata => i1137x_x2_2668,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2668
    phi_stmt_2674: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2677_wire & type_cast_2679_wire;
      req <= phi_stmt_2674_req_0 & phi_stmt_2674_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2674",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2674_ack_0,
          idata => idata,
          odata => j1187x_x1_2674,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2674
    phi_stmt_3001: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3004_wire & type_cast_3007_wire_constant;
      req <= phi_stmt_3001_req_0 & phi_stmt_3001_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3001",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3001_ack_0,
          idata => idata,
          odata => k1129x_x0x_xph_3001,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3001
    phi_stmt_3008: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3011_wire & type_cast_3013_wire;
      req <= phi_stmt_3008_req_0 & phi_stmt_3008_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3008",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3008_ack_0,
          idata => idata,
          odata => i1137x_x1x_xph_3008,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3008
    phi_stmt_3014: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3017_wire & type_cast_3019_wire;
      req <= phi_stmt_3014_req_0 & phi_stmt_3014_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3014",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3014_ack_0,
          idata => idata,
          odata => j1187x_x0x_xph_3014,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3014
    phi_stmt_3064: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3068_wire_constant & type_cast_3070_wire;
      req <= phi_stmt_3064_req_0 & phi_stmt_3064_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3064",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3064_ack_0,
          idata => idata,
          odata => k1351x_x1_3064,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3064
    phi_stmt_3071: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3074_wire & type_cast_3076_wire;
      req <= phi_stmt_3071_req_0 & phi_stmt_3071_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3071",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3071_ack_0,
          idata => idata,
          odata => i1355x_x2_3071,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3071
    phi_stmt_3077: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3080_wire & type_cast_3083_wire_constant;
      req <= phi_stmt_3077_req_0 & phi_stmt_3077_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3077",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3077_ack_0,
          idata => idata,
          odata => j1406x_x1_3077,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3077
    phi_stmt_338: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_342_wire_constant & type_cast_344_wire;
      req <= phi_stmt_338_req_0 & phi_stmt_338_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_338",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_338_ack_0,
          idata => idata,
          odata => indvar_338,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_338
    phi_stmt_3406: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3410_wire_constant & type_cast_3412_wire;
      req <= phi_stmt_3406_req_0 & phi_stmt_3406_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3406",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3406_ack_0,
          idata => idata,
          odata => k1351x_x0x_xph_3406,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3406
    phi_stmt_3413: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3416_wire & type_cast_3418_wire;
      req <= phi_stmt_3413_req_0 & phi_stmt_3413_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3413",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3413_ack_0,
          idata => idata,
          odata => i1355x_x1x_xph_3413,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3413
    phi_stmt_3419: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3422_wire & type_cast_3424_wire;
      req <= phi_stmt_3419_req_0 & phi_stmt_3419_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3419",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3419_ack_0,
          idata => idata,
          odata => j1406x_x0x_xph_3419,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3419
    phi_stmt_3475: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3479_wire_constant & type_cast_3481_wire;
      req <= phi_stmt_3475_req_0 & phi_stmt_3475_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3475",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3475_ack_0,
          idata => idata,
          odata => k1568x_x1_3475,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3475
    phi_stmt_3482: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3485_wire & type_cast_3487_wire;
      req <= phi_stmt_3482_req_0 & phi_stmt_3482_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3482",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3482_ack_0,
          idata => idata,
          odata => i1576x_x2_3482,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3482
    phi_stmt_3488: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3491_wire & type_cast_3493_wire;
      req <= phi_stmt_3488_req_0 & phi_stmt_3488_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3488",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3488_ack_0,
          idata => idata,
          odata => j1627x_x1_3488,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3488
    phi_stmt_3815: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3819_wire_constant & type_cast_3821_wire;
      req <= phi_stmt_3815_req_0 & phi_stmt_3815_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3815",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3815_ack_0,
          idata => idata,
          odata => k1568x_x0x_xph_3815,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3815
    phi_stmt_3822: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3825_wire & type_cast_3827_wire;
      req <= phi_stmt_3822_req_0 & phi_stmt_3822_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3822",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3822_ack_0,
          idata => idata,
          odata => i1576x_x1x_xph_3822,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3822
    phi_stmt_3828: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3831_wire & type_cast_3833_wire;
      req <= phi_stmt_3828_req_0 & phi_stmt_3828_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3828",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3828_ack_0,
          idata => idata,
          odata => j1627x_x0x_xph_3828,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3828
    phi_stmt_622: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_627_wire_constant & type_cast_629_wire;
      req <= phi_stmt_622_req_0 & phi_stmt_622_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_622",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_622_ack_0,
          idata => idata,
          odata => jx_x1_622,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_622
    phi_stmt_630: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_634_wire_constant & type_cast_636_wire;
      req <= phi_stmt_630_req_0 & phi_stmt_630_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_630",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_630_ack_0,
          idata => idata,
          odata => i68x_x2_630,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_630
    phi_stmt_637: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_641_wire_constant & type_cast_643_wire;
      req <= phi_stmt_637_req_0 & phi_stmt_637_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_637",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_637_ack_0,
          idata => idata,
          odata => kx_x1_637,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_637
    phi_stmt_967: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_970_wire & type_cast_972_wire;
      req <= phi_stmt_967_req_0 & phi_stmt_967_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_967",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_967_ack_0,
          idata => idata,
          odata => jx_x0x_xph_967,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_967
    phi_stmt_973: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_976_wire & type_cast_978_wire;
      req <= phi_stmt_973_req_0 & phi_stmt_973_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_973",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_973_ack_0,
          idata => idata,
          odata => i68x_x1x_xph_973,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_973
    phi_stmt_979: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_982_wire & type_cast_985_wire_constant;
      req <= phi_stmt_979_req_0 & phi_stmt_979_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_979",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_979_ack_0,
          idata => idata,
          odata => kx_x0x_xph_979,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_979
    -- flow-through select operator MUX_1356_inst
    j309x_x2_1357 <= div260_998 when (cmp443_1342(0) /=  '0') else inc434_1332;
    -- flow-through select operator MUX_1771_inst
    j525x_x2_1772 <= type_cast_1769_wire_constant when (cmp661_1756(0) /=  '0') else inc651_1746;
    -- flow-through select operator MUX_2168_inst
    j747x_x2_2169 <= div260_998 when (cmp881_2154(0) /=  '0') else inc872_2144;
    -- flow-through select operator MUX_2585_inst
    j963x_x2_2586 <= type_cast_2583_wire_constant when (cmp1100_2570(0) /=  '0') else inc1090_2560;
    -- flow-through select operator MUX_2982_inst
    j1187x_x2_2983 <= div260_998 when (cmp1322_2968(0) /=  '0') else inc1313_2958;
    -- flow-through select operator MUX_334_inst
    umax7_335 <= tmp5_322 when (tmp6_328(0) /=  '0') else type_cast_333_wire_constant;
    -- flow-through select operator MUX_3387_inst
    j1406x_x2_3388 <= type_cast_3385_wire_constant when (cmp1541_3372(0) /=  '0') else inc1531_3362;
    -- flow-through select operator MUX_3796_inst
    j1627x_x2_3797 <= div260_998 when (cmp1760_3782(0) /=  '0') else inc1751_3772;
    -- flow-through select operator MUX_948_inst
    jx_x2_949 <= type_cast_946_wire_constant when (cmp229_933(0) /=  '0') else inc219_923;
    addr_of_1178_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1178_final_reg_req_0;
      addr_of_1178_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1178_final_reg_req_1;
      addr_of_1178_final_reg_ack_1<= rack(0);
      addr_of_1178_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1178_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1177_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx368_1179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1261_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1261_final_reg_req_0;
      addr_of_1261_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1261_final_reg_req_1;
      addr_of_1261_final_reg_ack_1<= rack(0);
      addr_of_1261_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1261_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1260_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx411_1262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1286_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1286_final_reg_req_0;
      addr_of_1286_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1286_final_reg_req_1;
      addr_of_1286_final_reg_ack_1<= rack(0);
      addr_of_1286_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1286_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1285_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx416_1287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1592_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1592_final_reg_req_0;
      addr_of_1592_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1592_final_reg_req_1;
      addr_of_1592_final_reg_ack_1<= rack(0);
      addr_of_1592_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1592_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1591_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx585_1593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1675_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1675_final_reg_req_0;
      addr_of_1675_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1675_final_reg_req_1;
      addr_of_1675_final_reg_ack_1<= rack(0);
      addr_of_1675_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1675_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1674_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx628_1676,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1700_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1700_final_reg_req_0;
      addr_of_1700_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1700_final_reg_req_1;
      addr_of_1700_final_reg_ack_1<= rack(0);
      addr_of_1700_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1700_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1699_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx633_1701,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1990_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1990_final_reg_req_0;
      addr_of_1990_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1990_final_reg_req_1;
      addr_of_1990_final_reg_ack_1<= rack(0);
      addr_of_1990_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1990_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1989_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx806_1991,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2073_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2073_final_reg_req_0;
      addr_of_2073_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2073_final_reg_req_1;
      addr_of_2073_final_reg_ack_1<= rack(0);
      addr_of_2073_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2073_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2072_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx849_2074,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2098_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2098_final_reg_req_0;
      addr_of_2098_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2098_final_reg_req_1;
      addr_of_2098_final_reg_ack_1<= rack(0);
      addr_of_2098_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2098_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2097_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx854_2099,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2406_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2406_final_reg_req_0;
      addr_of_2406_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2406_final_reg_req_1;
      addr_of_2406_final_reg_ack_1<= rack(0);
      addr_of_2406_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2406_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2405_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1024_2407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2489_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2489_final_reg_req_0;
      addr_of_2489_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2489_final_reg_req_1;
      addr_of_2489_final_reg_ack_1<= rack(0);
      addr_of_2489_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2489_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2488_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1067_2490,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2514_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2514_final_reg_req_0;
      addr_of_2514_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2514_final_reg_req_1;
      addr_of_2514_final_reg_ack_1<= rack(0);
      addr_of_2514_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2514_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2513_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1072_2515,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2804_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2804_final_reg_req_0;
      addr_of_2804_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2804_final_reg_req_1;
      addr_of_2804_final_reg_ack_1<= rack(0);
      addr_of_2804_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2804_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2803_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1247_2805,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2887_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2887_final_reg_req_0;
      addr_of_2887_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2887_final_reg_req_1;
      addr_of_2887_final_reg_ack_1<= rack(0);
      addr_of_2887_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2887_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2886_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1290_2888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2912_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2912_final_reg_req_0;
      addr_of_2912_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2912_final_reg_req_1;
      addr_of_2912_final_reg_ack_1<= rack(0);
      addr_of_2912_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2912_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2911_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1295_2913,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3208_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3208_final_reg_req_0;
      addr_of_3208_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3208_final_reg_req_1;
      addr_of_3208_final_reg_ack_1<= rack(0);
      addr_of_3208_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3208_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3207_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1465_3209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3291_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3291_final_reg_req_0;
      addr_of_3291_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3291_final_reg_req_1;
      addr_of_3291_final_reg_ack_1<= rack(0);
      addr_of_3291_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3291_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3290_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1508_3292,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3316_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3316_final_reg_req_0;
      addr_of_3316_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3316_final_reg_req_1;
      addr_of_3316_final_reg_ack_1<= rack(0);
      addr_of_3316_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3316_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3315_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1513_3317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_351_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_351_final_reg_req_0;
      addr_of_351_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_351_final_reg_req_1;
      addr_of_351_final_reg_ack_1<= rack(0);
      addr_of_351_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_351_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_350_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3618_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3618_final_reg_req_0;
      addr_of_3618_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3618_final_reg_req_1;
      addr_of_3618_final_reg_ack_1<= rack(0);
      addr_of_3618_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3618_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3617_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1685_3619,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3701_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3701_final_reg_req_0;
      addr_of_3701_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3701_final_reg_req_1;
      addr_of_3701_final_reg_ack_1<= rack(0);
      addr_of_3701_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3701_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3700_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1728_3702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3726_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3726_final_reg_req_0;
      addr_of_3726_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3726_final_reg_req_1;
      addr_of_3726_final_reg_ack_1<= rack(0);
      addr_of_3726_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3726_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3725_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx1733_3727,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_769_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_769_final_reg_req_0;
      addr_of_769_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_769_final_reg_req_1;
      addr_of_769_final_reg_ack_1<= rack(0);
      addr_of_769_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_769_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_768_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx158_770,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_852_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_852_final_reg_req_0;
      addr_of_852_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_852_final_reg_req_1;
      addr_of_852_final_reg_ack_1<= rack(0);
      addr_of_852_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_852_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_851_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx198_853,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_877_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_877_final_reg_req_0;
      addr_of_877_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_877_final_reg_req_1;
      addr_of_877_final_reg_ack_1<= rack(0);
      addr_of_877_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_877_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_876_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx203_878,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1004_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1004_inst_req_0;
      type_cast_1004_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1004_inst_req_1;
      type_cast_1004_inst_ack_1<= rack(0);
      type_cast_1004_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1004_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp266_1001,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv317_1005,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1037_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1037_inst_req_0;
      type_cast_1037_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1037_inst_req_1;
      type_cast_1037_inst_ack_1<= rack(0);
      type_cast_1037_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1037_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div260_998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1037_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1039_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1039_inst_req_0;
      type_cast_1039_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1039_inst_req_1;
      type_cast_1039_inst_ack_1<= rack(0);
      type_cast_1039_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1039_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j309x_x0x_xph_1375,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1039_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1046_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1046_inst_req_0;
      type_cast_1046_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1046_inst_req_1;
      type_cast_1046_inst_ack_1<= rack(0);
      type_cast_1046_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1046_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i263x_x1x_xph_1381,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1046_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1053_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1053_inst_req_0;
      type_cast_1053_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1053_inst_req_1;
      type_cast_1053_inst_ack_1<= rack(0);
      type_cast_1053_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1053_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k255x_x0x_xph_1387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1053_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1058_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1058_inst_req_0;
      type_cast_1058_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1058_inst_req_1;
      type_cast_1058_inst_ack_1<= rack(0);
      type_cast_1058_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1058_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1057_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv315_1059,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1062_inst
    process(conv315_1059) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv315_1059(31 downto 0);
      type_cast_1062_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1064_inst
    process(conv317_1005) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv317_1005(31 downto 0);
      type_cast_1064_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1075_inst
    process(conv315_1059) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv315_1059(31 downto 0);
      type_cast_1075_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1077_inst
    process(add328_1026) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add328_1026(31 downto 0);
      type_cast_1077_wire <= tmp_var; -- 
    end process;
    type_cast_1095_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1095_inst_req_0;
      type_cast_1095_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1095_inst_req_1;
      type_cast_1095_inst_ack_1<= rack(0);
      type_cast_1095_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1095_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1094_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv333_1096,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1099_inst
    process(conv333_1096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv333_1096(31 downto 0);
      type_cast_1099_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1101_inst
    process(conv317_1005) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv317_1005(31 downto 0);
      type_cast_1101_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1112_inst
    process(conv333_1096) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv333_1096(31 downto 0);
      type_cast_1112_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1114_inst
    process(add345_1031) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add345_1031(31 downto 0);
      type_cast_1114_wire <= tmp_var; -- 
    end process;
    type_cast_1132_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1132_inst_req_0;
      type_cast_1132_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1132_inst_req_1;
      type_cast_1132_inst_ack_1<= rack(0);
      type_cast_1132_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1132_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1131_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv352_1133,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1137_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1137_inst_req_0;
      type_cast_1137_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1137_inst_req_1;
      type_cast_1137_inst_ack_1<= rack(0);
      type_cast_1137_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1137_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1136_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv356_1138,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1161_inst
    process(add364_1158) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add364_1158(31 downto 0);
      type_cast_1161_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1166_inst
    process(ASHR_i32_i32_1165_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1165_wire(31 downto 0);
      shr366_1167 <= tmp_var; -- 
    end process;
    type_cast_1171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1171_inst_req_0;
      type_cast_1171_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1171_inst_req_1;
      type_cast_1171_inst_ack_1<= rack(0);
      type_cast_1171_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1171_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1170_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom367_1172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1190_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1190_inst_req_0;
      type_cast_1190_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1190_inst_req_1;
      type_cast_1190_inst_ack_1<= rack(0);
      type_cast_1190_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1190_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1189_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv373_1191,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1244_inst
    process(add391_1221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add391_1221(31 downto 0);
      type_cast_1244_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1249_inst
    process(ASHR_i32_i32_1248_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1248_wire(31 downto 0);
      shr409_1250 <= tmp_var; -- 
    end process;
    type_cast_1254_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1254_inst_req_0;
      type_cast_1254_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1254_inst_req_1;
      type_cast_1254_inst_ack_1<= rack(0);
      type_cast_1254_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1254_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1253_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom410_1255,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1269_inst
    process(add407_1241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add407_1241(31 downto 0);
      type_cast_1269_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1274_inst
    process(ASHR_i32_i32_1273_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1273_wire(31 downto 0);
      shr414_1275 <= tmp_var; -- 
    end process;
    type_cast_1279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1279_inst_req_0;
      type_cast_1279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1279_inst_req_1;
      type_cast_1279_inst_ack_1<= rack(0);
      type_cast_1279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1278_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom415_1280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1297_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1297_inst_req_0;
      type_cast_1297_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1297_inst_req_1;
      type_cast_1297_inst_ack_1<= rack(0);
      type_cast_1297_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1297_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1296_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv421_1298,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1307_inst
    process(add422_1304) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add422_1304(31 downto 0);
      type_cast_1307_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1309_inst
    process(conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv92_517(31 downto 0);
      type_cast_1309_wire <= tmp_var; -- 
    end process;
    type_cast_1336_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1336_inst_req_0;
      type_cast_1336_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1336_inst_req_1;
      type_cast_1336_inst_ack_1<= rack(0);
      type_cast_1336_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1336_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1335_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv436_1337,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1345_inst_req_0;
      type_cast_1345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1345_inst_req_1;
      type_cast_1345_inst_ack_1<= rack(0);
      type_cast_1345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp443_1342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc448_1346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1361_inst_req_0;
      type_cast_1361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1361_inst_req_1;
      type_cast_1361_inst_ack_1<= rack(0);
      type_cast_1361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1360_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv451_1362,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1378_inst_req_0;
      type_cast_1378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1378_inst_req_1;
      type_cast_1378_inst_ack_1<= rack(0);
      type_cast_1378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j309x_x1_1034,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1378_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1380_inst_req_0;
      type_cast_1380_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1380_inst_req_1;
      type_cast_1380_inst_ack_1<= rack(0);
      type_cast_1380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j309x_x2_1357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1380_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1384_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1384_inst_req_0;
      type_cast_1384_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1384_inst_req_1;
      type_cast_1384_inst_ack_1<= rack(0);
      type_cast_1384_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1384_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i263x_x2_1040,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1384_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1386_inst_req_0;
      type_cast_1386_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1386_inst_req_1;
      type_cast_1386_inst_ack_1<= rack(0);
      type_cast_1386_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc448x_xi263x_x2_1351,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1386_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1390_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1390_inst_req_0;
      type_cast_1390_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1390_inst_req_1;
      type_cast_1390_inst_ack_1<= rack(0);
      type_cast_1390_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1390_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add430_1324,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1390_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1399_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1399_inst_req_0;
      type_cast_1399_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1399_inst_req_1;
      type_cast_1399_inst_ack_1<= rack(0);
      type_cast_1399_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1399_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv477_1400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1412_inst_req_0;
      type_cast_1412_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1412_inst_req_1;
      type_cast_1412_inst_ack_1<= rack(0);
      type_cast_1412_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1412_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp482_1409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv533_1413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1454_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1454_inst_req_0;
      type_cast_1454_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1454_inst_req_1;
      type_cast_1454_inst_ack_1<= rack(0);
      type_cast_1454_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1454_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k471x_x0x_xph_1790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1454_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1458_inst_req_0;
      type_cast_1458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1458_inst_req_1;
      type_cast_1458_inst_ack_1<= rack(0);
      type_cast_1458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1458_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div478_1406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1458_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1460_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1460_inst_req_0;
      type_cast_1460_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1460_inst_req_1;
      type_cast_1460_inst_ack_1<= rack(0);
      type_cast_1460_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1460_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i475x_x1x_xph_1797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1460_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1467_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1467_inst_req_0;
      type_cast_1467_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1467_inst_req_1;
      type_cast_1467_inst_ack_1<= rack(0);
      type_cast_1467_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1467_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j525x_x0x_xph_1803,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1467_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1472_inst_req_0;
      type_cast_1472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1472_inst_req_1;
      type_cast_1472_inst_ack_1<= rack(0);
      type_cast_1472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1471_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv531_1473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1476_inst
    process(conv531_1473) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv531_1473(31 downto 0);
      type_cast_1476_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1478_inst
    process(conv533_1413) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv533_1413(31 downto 0);
      type_cast_1478_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1489_inst
    process(conv531_1473) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv531_1473(31 downto 0);
      type_cast_1489_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1491_inst
    process(add544_1440) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add544_1440(31 downto 0);
      type_cast_1491_wire <= tmp_var; -- 
    end process;
    type_cast_1509_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1509_inst_req_0;
      type_cast_1509_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1509_inst_req_1;
      type_cast_1509_inst_ack_1<= rack(0);
      type_cast_1509_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1509_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1508_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv549_1510,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1513_inst
    process(conv549_1510) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv549_1510(31 downto 0);
      type_cast_1513_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1515_inst
    process(conv533_1413) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv533_1413(31 downto 0);
      type_cast_1515_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1526_inst
    process(conv549_1510) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv549_1510(31 downto 0);
      type_cast_1526_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1528_inst
    process(add562_1445) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add562_1445(31 downto 0);
      type_cast_1528_wire <= tmp_var; -- 
    end process;
    type_cast_1546_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1546_inst_req_0;
      type_cast_1546_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1546_inst_req_1;
      type_cast_1546_inst_ack_1<= rack(0);
      type_cast_1546_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1546_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1545_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv569_1547,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1551_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1551_inst_req_0;
      type_cast_1551_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1551_inst_req_1;
      type_cast_1551_inst_ack_1<= rack(0);
      type_cast_1551_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1551_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1550_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv573_1552,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1575_inst
    process(add581_1572) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add581_1572(31 downto 0);
      type_cast_1575_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1580_inst
    process(ASHR_i32_i32_1579_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1579_wire(31 downto 0);
      shr583_1581 <= tmp_var; -- 
    end process;
    type_cast_1585_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1585_inst_req_0;
      type_cast_1585_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1585_inst_req_1;
      type_cast_1585_inst_ack_1<= rack(0);
      type_cast_1585_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1585_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1584_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom584_1586,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1604_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1604_inst_req_0;
      type_cast_1604_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1604_inst_req_1;
      type_cast_1604_inst_ack_1<= rack(0);
      type_cast_1604_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1604_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1603_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv590_1605,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1658_inst
    process(add608_1635) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add608_1635(31 downto 0);
      type_cast_1658_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1663_inst
    process(ASHR_i32_i32_1662_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1662_wire(31 downto 0);
      shr626_1664 <= tmp_var; -- 
    end process;
    type_cast_1668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1668_inst_req_0;
      type_cast_1668_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1668_inst_req_1;
      type_cast_1668_inst_ack_1<= rack(0);
      type_cast_1668_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1668_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1667_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom627_1669,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1683_inst
    process(add624_1655) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add624_1655(31 downto 0);
      type_cast_1683_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1688_inst
    process(ASHR_i32_i32_1687_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1687_wire(31 downto 0);
      shr631_1689 <= tmp_var; -- 
    end process;
    type_cast_1693_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1693_inst_req_0;
      type_cast_1693_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1693_inst_req_1;
      type_cast_1693_inst_ack_1<= rack(0);
      type_cast_1693_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1693_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1692_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom632_1694,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1711_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1711_inst_req_0;
      type_cast_1711_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1711_inst_req_1;
      type_cast_1711_inst_ack_1<= rack(0);
      type_cast_1711_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1711_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1710_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv638_1712,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1721_inst
    process(add639_1718) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add639_1718(31 downto 0);
      type_cast_1721_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1723_inst
    process(conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv92_517(31 downto 0);
      type_cast_1723_wire <= tmp_var; -- 
    end process;
    type_cast_1750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1750_inst_req_0;
      type_cast_1750_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1750_inst_req_1;
      type_cast_1750_inst_ack_1<= rack(0);
      type_cast_1750_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1750_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1749_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv653_1751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1759_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1759_inst_req_0;
      type_cast_1759_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1759_inst_req_1;
      type_cast_1759_inst_ack_1<= rack(0);
      type_cast_1759_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1759_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp661_1756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc666_1760,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1776_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1776_inst_req_0;
      type_cast_1776_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1776_inst_req_1;
      type_cast_1776_inst_ack_1<= rack(0);
      type_cast_1776_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1776_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1775_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv669_1777,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1793_inst_req_0;
      type_cast_1793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1793_inst_req_1;
      type_cast_1793_inst_ack_1<= rack(0);
      type_cast_1793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add647_1738,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1793_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1800_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1800_inst_req_0;
      type_cast_1800_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1800_inst_req_1;
      type_cast_1800_inst_ack_1<= rack(0);
      type_cast_1800_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1800_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i475x_x2_1455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1800_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1802_inst_req_0;
      type_cast_1802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1802_inst_req_1;
      type_cast_1802_inst_ack_1<= rack(0);
      type_cast_1802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc666x_xi475x_x2_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1802_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1806_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1806_inst_req_0;
      type_cast_1806_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1806_inst_req_1;
      type_cast_1806_inst_ack_1<= rack(0);
      type_cast_1806_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1806_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j525x_x1_1461,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1806_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1808_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1808_inst_req_0;
      type_cast_1808_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1808_inst_req_1;
      type_cast_1808_inst_ack_1<= rack(0);
      type_cast_1808_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1808_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j525x_x2_1772,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1808_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1817_inst_req_0;
      type_cast_1817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1817_inst_req_1;
      type_cast_1817_inst_ack_1<= rack(0);
      type_cast_1817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp704_1814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv755_1818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1850_inst_req_0;
      type_cast_1850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1850_inst_req_1;
      type_cast_1850_inst_ack_1<= rack(0);
      type_cast_1850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k689x_x0x_xph_2187,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1850_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1857_inst_req_0;
      type_cast_1857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1857_inst_req_1;
      type_cast_1857_inst_ack_1<= rack(0);
      type_cast_1857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i697x_x1x_xph_2194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1857_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1859_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1859_inst_req_0;
      type_cast_1859_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1859_inst_req_1;
      type_cast_1859_inst_ack_1<= rack(0);
      type_cast_1859_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1859_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div478_1406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1859_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1863_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1863_inst_req_0;
      type_cast_1863_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1863_inst_req_1;
      type_cast_1863_inst_ack_1<= rack(0);
      type_cast_1863_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1863_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j747x_x0x_xph_2200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1863_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1865_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1865_inst_req_0;
      type_cast_1865_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1865_inst_req_1;
      type_cast_1865_inst_ack_1<= rack(0);
      type_cast_1865_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1865_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div260_998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1865_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1870_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1870_inst_req_0;
      type_cast_1870_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1870_inst_req_1;
      type_cast_1870_inst_ack_1<= rack(0);
      type_cast_1870_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1870_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1869_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv753_1871,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1874_inst
    process(conv753_1871) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv753_1871(31 downto 0);
      type_cast_1874_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1876_inst
    process(conv755_1818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv755_1818(31 downto 0);
      type_cast_1876_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1887_inst
    process(conv753_1871) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv753_1871(31 downto 0);
      type_cast_1887_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1889_inst
    process(add766_1839) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add766_1839(31 downto 0);
      type_cast_1889_wire <= tmp_var; -- 
    end process;
    type_cast_1907_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1907_inst_req_0;
      type_cast_1907_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1907_inst_req_1;
      type_cast_1907_inst_ack_1<= rack(0);
      type_cast_1907_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1907_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1906_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv771_1908,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1911_inst
    process(conv771_1908) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv771_1908(31 downto 0);
      type_cast_1911_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1913_inst
    process(conv755_1818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv755_1818(31 downto 0);
      type_cast_1913_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1924_inst
    process(conv771_1908) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv771_1908(31 downto 0);
      type_cast_1924_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1926_inst
    process(add783_1844) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add783_1844(31 downto 0);
      type_cast_1926_wire <= tmp_var; -- 
    end process;
    type_cast_1944_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1944_inst_req_0;
      type_cast_1944_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1944_inst_req_1;
      type_cast_1944_inst_ack_1<= rack(0);
      type_cast_1944_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1944_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1943_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv790_1945,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1949_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1949_inst_req_0;
      type_cast_1949_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1949_inst_req_1;
      type_cast_1949_inst_ack_1<= rack(0);
      type_cast_1949_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1949_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1948_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv794_1950,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1973_inst
    process(add802_1970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add802_1970(31 downto 0);
      type_cast_1973_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1978_inst
    process(ASHR_i32_i32_1977_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1977_wire(31 downto 0);
      shr804_1979 <= tmp_var; -- 
    end process;
    type_cast_1983_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1983_inst_req_0;
      type_cast_1983_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1983_inst_req_1;
      type_cast_1983_inst_ack_1<= rack(0);
      type_cast_1983_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1983_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1982_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom805_1984,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2002_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2002_inst_req_0;
      type_cast_2002_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2002_inst_req_1;
      type_cast_2002_inst_ack_1<= rack(0);
      type_cast_2002_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2002_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2001_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv811_2003,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2056_inst
    process(add829_2033) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add829_2033(31 downto 0);
      type_cast_2056_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2061_inst
    process(ASHR_i32_i32_2060_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2060_wire(31 downto 0);
      shr847_2062 <= tmp_var; -- 
    end process;
    type_cast_2066_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2066_inst_req_0;
      type_cast_2066_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2066_inst_req_1;
      type_cast_2066_inst_ack_1<= rack(0);
      type_cast_2066_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2066_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2065_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom848_2067,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2081_inst
    process(add845_2053) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add845_2053(31 downto 0);
      type_cast_2081_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2086_inst
    process(ASHR_i32_i32_2085_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2085_wire(31 downto 0);
      shr852_2087 <= tmp_var; -- 
    end process;
    type_cast_2091_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2091_inst_req_0;
      type_cast_2091_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2091_inst_req_1;
      type_cast_2091_inst_ack_1<= rack(0);
      type_cast_2091_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2091_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2090_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom853_2092,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2109_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2109_inst_req_0;
      type_cast_2109_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2109_inst_req_1;
      type_cast_2109_inst_ack_1<= rack(0);
      type_cast_2109_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2109_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2108_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv859_2110,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2119_inst
    process(add860_2116) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add860_2116(31 downto 0);
      type_cast_2119_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2121_inst
    process(conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv92_517(31 downto 0);
      type_cast_2121_wire <= tmp_var; -- 
    end process;
    type_cast_2148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2148_inst_req_0;
      type_cast_2148_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2148_inst_req_1;
      type_cast_2148_inst_ack_1<= rack(0);
      type_cast_2148_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2148_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2147_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv874_2149,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2157_inst_req_0;
      type_cast_2157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2157_inst_req_1;
      type_cast_2157_inst_ack_1<= rack(0);
      type_cast_2157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp881_2154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc886_2158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2173_inst_req_0;
      type_cast_2173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2173_inst_req_1;
      type_cast_2173_inst_ack_1<= rack(0);
      type_cast_2173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2172_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv889_2174,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2193_inst_req_0;
      type_cast_2193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2193_inst_req_1;
      type_cast_2193_inst_ack_1<= rack(0);
      type_cast_2193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add868_2136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2193_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2197_inst_req_0;
      type_cast_2197_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2197_inst_req_1;
      type_cast_2197_inst_ack_1<= rack(0);
      type_cast_2197_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2197_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i697x_x2_1854,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2197_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2199_inst_req_0;
      type_cast_2199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2199_inst_req_1;
      type_cast_2199_inst_ack_1<= rack(0);
      type_cast_2199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc886x_xi697x_x2_2163,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2199_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2203_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2203_inst_req_0;
      type_cast_2203_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2203_inst_req_1;
      type_cast_2203_inst_ack_1<= rack(0);
      type_cast_2203_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2203_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j747x_x2_2169,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2203_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2205_inst_req_0;
      type_cast_2205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2205_inst_req_1;
      type_cast_2205_inst_ack_1<= rack(0);
      type_cast_2205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j747x_x1_1860,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2205_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2220_inst_req_0;
      type_cast_2220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2220_inst_req_1;
      type_cast_2220_inst_ack_1<= rack(0);
      type_cast_2220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp920_2217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv971_2221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2268_inst_req_0;
      type_cast_2268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2268_inst_req_1;
      type_cast_2268_inst_ack_1<= rack(0);
      type_cast_2268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k909x_x0x_xph_2604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2268_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2272_inst_req_0;
      type_cast_2272_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2272_inst_req_1;
      type_cast_2272_inst_ack_1<= rack(0);
      type_cast_2272_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2272_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div916_2214,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2272_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2274_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2274_inst_req_0;
      type_cast_2274_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2274_inst_req_1;
      type_cast_2274_inst_ack_1<= rack(0);
      type_cast_2274_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2274_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i913x_x1x_xph_2611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2274_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2281_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2281_inst_req_0;
      type_cast_2281_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2281_inst_req_1;
      type_cast_2281_inst_ack_1<= rack(0);
      type_cast_2281_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2281_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j963x_x0x_xph_2617,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2281_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2286_inst_req_0;
      type_cast_2286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2286_inst_req_1;
      type_cast_2286_inst_ack_1<= rack(0);
      type_cast_2286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2285_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv969_2287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2290_inst
    process(conv969_2287) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv969_2287(31 downto 0);
      type_cast_2290_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2292_inst
    process(conv971_2221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv971_2221(31 downto 0);
      type_cast_2292_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2303_inst
    process(conv969_2287) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv969_2287(31 downto 0);
      type_cast_2303_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2305_inst
    process(add983_2254) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add983_2254(31 downto 0);
      type_cast_2305_wire <= tmp_var; -- 
    end process;
    type_cast_2323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2323_inst_req_0;
      type_cast_2323_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2323_inst_req_1;
      type_cast_2323_inst_ack_1<= rack(0);
      type_cast_2323_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2323_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2322_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv988_2324,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2327_inst
    process(conv988_2324) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv988_2324(31 downto 0);
      type_cast_2327_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2329_inst
    process(conv971_2221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv971_2221(31 downto 0);
      type_cast_2329_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2340_inst
    process(conv988_2324) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv988_2324(31 downto 0);
      type_cast_2340_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2342_inst
    process(add1001_2259) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1001_2259(31 downto 0);
      type_cast_2342_wire <= tmp_var; -- 
    end process;
    type_cast_2360_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2360_inst_req_0;
      type_cast_2360_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2360_inst_req_1;
      type_cast_2360_inst_ack_1<= rack(0);
      type_cast_2360_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2360_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2359_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1008_2361,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2365_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2365_inst_req_0;
      type_cast_2365_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2365_inst_req_1;
      type_cast_2365_inst_ack_1<= rack(0);
      type_cast_2365_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2365_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2364_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1012_2366,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2389_inst
    process(add1020_2386) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1020_2386(31 downto 0);
      type_cast_2389_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2394_inst
    process(ASHR_i32_i32_2393_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2393_wire(31 downto 0);
      shr1022_2395 <= tmp_var; -- 
    end process;
    type_cast_2399_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2399_inst_req_0;
      type_cast_2399_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2399_inst_req_1;
      type_cast_2399_inst_ack_1<= rack(0);
      type_cast_2399_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2399_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2398_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1023_2400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2418_inst_req_0;
      type_cast_2418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2418_inst_req_1;
      type_cast_2418_inst_ack_1<= rack(0);
      type_cast_2418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2417_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1029_2419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2472_inst
    process(add1047_2449) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1047_2449(31 downto 0);
      type_cast_2472_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2477_inst
    process(ASHR_i32_i32_2476_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2476_wire(31 downto 0);
      shr1065_2478 <= tmp_var; -- 
    end process;
    type_cast_2482_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2482_inst_req_0;
      type_cast_2482_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2482_inst_req_1;
      type_cast_2482_inst_ack_1<= rack(0);
      type_cast_2482_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2482_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2481_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1066_2483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2497_inst
    process(add1063_2469) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1063_2469(31 downto 0);
      type_cast_2497_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2502_inst
    process(ASHR_i32_i32_2501_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2501_wire(31 downto 0);
      shr1070_2503 <= tmp_var; -- 
    end process;
    type_cast_2507_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2507_inst_req_0;
      type_cast_2507_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2507_inst_req_1;
      type_cast_2507_inst_ack_1<= rack(0);
      type_cast_2507_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2507_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2506_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1071_2508,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2525_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2525_inst_req_0;
      type_cast_2525_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2525_inst_req_1;
      type_cast_2525_inst_ack_1<= rack(0);
      type_cast_2525_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2525_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2524_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1077_2526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2535_inst
    process(add1078_2532) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1078_2532(31 downto 0);
      type_cast_2535_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2537_inst
    process(conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv92_517(31 downto 0);
      type_cast_2537_wire <= tmp_var; -- 
    end process;
    type_cast_2564_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2564_inst_req_0;
      type_cast_2564_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2564_inst_req_1;
      type_cast_2564_inst_ack_1<= rack(0);
      type_cast_2564_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2564_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2563_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1092_2565,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_256_inst_req_0;
      type_cast_256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_256_inst_req_1;
      type_cast_256_inst_ack_1<= rack(0);
      type_cast_256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2573_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2573_inst_req_0;
      type_cast_2573_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2573_inst_req_1;
      type_cast_2573_inst_ack_1<= rack(0);
      type_cast_2573_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2573_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1100_2570,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1105_2574,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2590_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2590_inst_req_0;
      type_cast_2590_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2590_inst_req_1;
      type_cast_2590_inst_ack_1<= rack(0);
      type_cast_2590_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2590_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2589_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1108_2591,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2607_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2607_inst_req_0;
      type_cast_2607_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2607_inst_req_1;
      type_cast_2607_inst_ack_1<= rack(0);
      type_cast_2607_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2607_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1086_2552,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2607_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_260_inst_req_0;
      type_cast_260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_260_inst_req_1;
      type_cast_260_inst_ack_1<= rack(0);
      type_cast_260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10_261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2614_inst_req_0;
      type_cast_2614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2614_inst_req_1;
      type_cast_2614_inst_ack_1<= rack(0);
      type_cast_2614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i913x_x2_2269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2614_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2616_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2616_inst_req_0;
      type_cast_2616_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2616_inst_req_1;
      type_cast_2616_inst_ack_1<= rack(0);
      type_cast_2616_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2616_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1105x_xi913x_x2_2579,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2616_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2620_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2620_inst_req_0;
      type_cast_2620_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2620_inst_req_1;
      type_cast_2620_inst_ack_1<= rack(0);
      type_cast_2620_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2620_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j963x_x1_2275,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2620_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2622_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2622_inst_req_0;
      type_cast_2622_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2622_inst_req_1;
      type_cast_2622_inst_ack_1<= rack(0);
      type_cast_2622_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2622_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j963x_x2_2586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2622_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2631_inst_req_0;
      type_cast_2631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2631_inst_req_1;
      type_cast_2631_inst_ack_1<= rack(0);
      type_cast_2631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1144_2628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1195_2632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_264_inst_req_0;
      type_cast_264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_264_inst_req_1;
      type_cast_264_inst_ack_1<= rack(0);
      type_cast_264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_264_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_265,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2667_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2667_inst_req_0;
      type_cast_2667_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2667_inst_req_1;
      type_cast_2667_inst_ack_1<= rack(0);
      type_cast_2667_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2667_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1129x_x0x_xph_3001,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2667_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2671_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2671_inst_req_0;
      type_cast_2671_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2671_inst_req_1;
      type_cast_2671_inst_ack_1<= rack(0);
      type_cast_2671_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2671_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div916_2214,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2671_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2673_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2673_inst_req_0;
      type_cast_2673_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2673_inst_req_1;
      type_cast_2673_inst_ack_1<= rack(0);
      type_cast_2673_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2673_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1137x_x1x_xph_3008,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2673_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2677_inst_req_0;
      type_cast_2677_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2677_inst_req_1;
      type_cast_2677_inst_ack_1<= rack(0);
      type_cast_2677_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2677_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div260_998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2677_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2679_inst_req_0;
      type_cast_2679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2679_inst_req_1;
      type_cast_2679_inst_ack_1<= rack(0);
      type_cast_2679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2679_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1187x_x0x_xph_3014,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2679_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2684_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2684_inst_req_0;
      type_cast_2684_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2684_inst_req_1;
      type_cast_2684_inst_ack_1<= rack(0);
      type_cast_2684_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2684_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2683_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1193_2685,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2688_inst
    process(conv1193_2685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1193_2685(31 downto 0);
      type_cast_2688_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2690_inst
    process(conv1195_2632) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1195_2632(31 downto 0);
      type_cast_2690_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2701_inst
    process(conv1193_2685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1193_2685(31 downto 0);
      type_cast_2701_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2703_inst
    process(add1207_2653) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1207_2653(31 downto 0);
      type_cast_2703_wire <= tmp_var; -- 
    end process;
    type_cast_2721_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2721_inst_req_0;
      type_cast_2721_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2721_inst_req_1;
      type_cast_2721_inst_ack_1<= rack(0);
      type_cast_2721_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2721_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2720_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1212_2722,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2725_inst
    process(conv1212_2722) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1212_2722(31 downto 0);
      type_cast_2725_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2727_inst
    process(conv1195_2632) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1195_2632(31 downto 0);
      type_cast_2727_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2738_inst
    process(conv1212_2722) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1212_2722(31 downto 0);
      type_cast_2738_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2740_inst
    process(add1224_2658) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1224_2658(31 downto 0);
      type_cast_2740_wire <= tmp_var; -- 
    end process;
    type_cast_2758_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2758_inst_req_0;
      type_cast_2758_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2758_inst_req_1;
      type_cast_2758_inst_ack_1<= rack(0);
      type_cast_2758_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2758_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2757_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1231_2759,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2763_inst_req_0;
      type_cast_2763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2763_inst_req_1;
      type_cast_2763_inst_ack_1<= rack(0);
      type_cast_2763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2762_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1235_2764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2787_inst
    process(add1243_2784) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1243_2784(31 downto 0);
      type_cast_2787_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2792_inst
    process(ASHR_i32_i32_2791_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2791_wire(31 downto 0);
      shr1245_2793 <= tmp_var; -- 
    end process;
    type_cast_2797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2797_inst_req_0;
      type_cast_2797_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2797_inst_req_1;
      type_cast_2797_inst_ack_1<= rack(0);
      type_cast_2797_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2797_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2796_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1246_2798,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2816_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2816_inst_req_0;
      type_cast_2816_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2816_inst_req_1;
      type_cast_2816_inst_ack_1<= rack(0);
      type_cast_2816_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2816_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2815_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1252_2817,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2870_inst
    process(add1270_2847) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1270_2847(31 downto 0);
      type_cast_2870_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2875_inst
    process(ASHR_i32_i32_2874_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2874_wire(31 downto 0);
      shr1288_2876 <= tmp_var; -- 
    end process;
    type_cast_2880_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2880_inst_req_0;
      type_cast_2880_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2880_inst_req_1;
      type_cast_2880_inst_ack_1<= rack(0);
      type_cast_2880_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2880_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2879_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1289_2881,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2895_inst
    process(add1286_2867) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1286_2867(31 downto 0);
      type_cast_2895_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2900_inst
    process(ASHR_i32_i32_2899_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2899_wire(31 downto 0);
      shr1293_2901 <= tmp_var; -- 
    end process;
    type_cast_2905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2905_inst_req_0;
      type_cast_2905_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2905_inst_req_1;
      type_cast_2905_inst_ack_1<= rack(0);
      type_cast_2905_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2905_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2904_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1294_2906,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2923_inst_req_0;
      type_cast_2923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2923_inst_req_1;
      type_cast_2923_inst_ack_1<= rack(0);
      type_cast_2923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2922_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1300_2924,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2933_inst
    process(add1301_2930) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1301_2930(31 downto 0);
      type_cast_2933_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2935_inst
    process(conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv92_517(31 downto 0);
      type_cast_2935_wire <= tmp_var; -- 
    end process;
    type_cast_2962_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2962_inst_req_0;
      type_cast_2962_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2962_inst_req_1;
      type_cast_2962_inst_ack_1<= rack(0);
      type_cast_2962_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2962_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2961_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1315_2963,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2971_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2971_inst_req_0;
      type_cast_2971_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2971_inst_req_1;
      type_cast_2971_inst_ack_1<= rack(0);
      type_cast_2971_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2971_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1322_2968,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1327_2972,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_297_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_297_inst_req_0;
      type_cast_297_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_297_inst_req_1;
      type_cast_297_inst_ack_1<= rack(0);
      type_cast_297_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_297_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp_298,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2987_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2987_inst_req_0;
      type_cast_2987_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2987_inst_req_1;
      type_cast_2987_inst_ack_1<= rack(0);
      type_cast_2987_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2987_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2986_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1330_2988,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3004_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3004_inst_req_0;
      type_cast_3004_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3004_inst_req_1;
      type_cast_3004_inst_ack_1<= rack(0);
      type_cast_3004_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3004_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1309_2950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3004_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3011_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3011_inst_req_0;
      type_cast_3011_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3011_inst_req_1;
      type_cast_3011_inst_ack_1<= rack(0);
      type_cast_3011_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3011_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1137x_x2_2668,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3011_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3013_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3013_inst_req_0;
      type_cast_3013_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3013_inst_req_1;
      type_cast_3013_inst_ack_1<= rack(0);
      type_cast_3013_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3013_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1327x_xi1137x_x2_2977,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3013_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3017_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3017_inst_req_0;
      type_cast_3017_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3017_inst_req_1;
      type_cast_3017_inst_ack_1<= rack(0);
      type_cast_3017_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3017_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1187x_x1_2674,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3017_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3019_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3019_inst_req_0;
      type_cast_3019_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3019_inst_req_1;
      type_cast_3019_inst_ack_1<= rack(0);
      type_cast_3019_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3019_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1187x_x2_2983,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3019_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_301_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_301_inst_req_0;
      type_cast_301_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_301_inst_req_1;
      type_cast_301_inst_ack_1<= rack(0);
      type_cast_301_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_301_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_302,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3034_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3034_inst_req_0;
      type_cast_3034_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3034_inst_req_1;
      type_cast_3034_inst_ack_1<= rack(0);
      type_cast_3034_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3034_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1363_3031,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1414_3035,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3070_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3070_inst_req_0;
      type_cast_3070_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3070_inst_req_1;
      type_cast_3070_inst_ack_1<= rack(0);
      type_cast_3070_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3070_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1351x_x0x_xph_3406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3070_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3074_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3074_inst_req_0;
      type_cast_3074_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3074_inst_req_1;
      type_cast_3074_inst_ack_1<= rack(0);
      type_cast_3074_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3074_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1355x_x1x_xph_3413,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3074_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3076_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3076_inst_req_0;
      type_cast_3076_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3076_inst_req_1;
      type_cast_3076_inst_ack_1<= rack(0);
      type_cast_3076_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3076_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul1359_3028,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3076_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3080_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3080_inst_req_0;
      type_cast_3080_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3080_inst_req_1;
      type_cast_3080_inst_ack_1<= rack(0);
      type_cast_3080_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3080_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1406x_x0x_xph_3419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3080_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3088_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3088_inst_req_0;
      type_cast_3088_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3088_inst_req_1;
      type_cast_3088_inst_ack_1<= rack(0);
      type_cast_3088_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3088_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3087_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1412_3089,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3092_inst
    process(conv1412_3089) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1412_3089(31 downto 0);
      type_cast_3092_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3094_inst
    process(conv1414_3035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1414_3035(31 downto 0);
      type_cast_3094_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3105_inst
    process(conv1412_3089) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1412_3089(31 downto 0);
      type_cast_3105_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3107_inst
    process(add1424_3056) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1424_3056(31 downto 0);
      type_cast_3107_wire <= tmp_var; -- 
    end process;
    type_cast_310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_310_inst_req_0;
      type_cast_310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_310_inst_req_1;
      type_cast_310_inst_ack_1<= rack(0);
      type_cast_310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3125_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3125_inst_req_0;
      type_cast_3125_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3125_inst_req_1;
      type_cast_3125_inst_ack_1<= rack(0);
      type_cast_3125_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3125_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3124_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1429_3126,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3129_inst
    process(conv1429_3126) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1429_3126(31 downto 0);
      type_cast_3129_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3131_inst
    process(conv1414_3035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1414_3035(31 downto 0);
      type_cast_3131_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3142_inst
    process(conv1429_3126) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1429_3126(31 downto 0);
      type_cast_3142_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3144_inst
    process(add1442_3061) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1442_3061(31 downto 0);
      type_cast_3144_wire <= tmp_var; -- 
    end process;
    type_cast_3162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3162_inst_req_0;
      type_cast_3162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3162_inst_req_1;
      type_cast_3162_inst_ack_1<= rack(0);
      type_cast_3162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3161_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1449_3163,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3167_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3167_inst_req_0;
      type_cast_3167_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3167_inst_req_1;
      type_cast_3167_inst_ack_1<= rack(0);
      type_cast_3167_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3167_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3166_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1453_3168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3191_inst
    process(add1461_3188) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1461_3188(31 downto 0);
      type_cast_3191_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3196_inst
    process(ASHR_i32_i32_3195_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3195_wire(31 downto 0);
      shr1463_3197 <= tmp_var; -- 
    end process;
    type_cast_3201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3201_inst_req_0;
      type_cast_3201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3201_inst_req_1;
      type_cast_3201_inst_ack_1<= rack(0);
      type_cast_3201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3200_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1464_3202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3220_inst_req_0;
      type_cast_3220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3220_inst_req_1;
      type_cast_3220_inst_ack_1<= rack(0);
      type_cast_3220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3219_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1470_3221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3274_inst
    process(add1488_3251) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1488_3251(31 downto 0);
      type_cast_3274_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3279_inst
    process(ASHR_i32_i32_3278_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3278_wire(31 downto 0);
      shr1506_3280 <= tmp_var; -- 
    end process;
    type_cast_3284_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3284_inst_req_0;
      type_cast_3284_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3284_inst_req_1;
      type_cast_3284_inst_ack_1<= rack(0);
      type_cast_3284_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3284_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3283_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1507_3285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3299_inst
    process(add1504_3271) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1504_3271(31 downto 0);
      type_cast_3299_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3304_inst
    process(ASHR_i32_i32_3303_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3303_wire(31 downto 0);
      shr1511_3305 <= tmp_var; -- 
    end process;
    type_cast_3309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3309_inst_req_0;
      type_cast_3309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3309_inst_req_1;
      type_cast_3309_inst_ack_1<= rack(0);
      type_cast_3309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3308_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1512_3310,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3327_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3327_inst_req_0;
      type_cast_3327_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3327_inst_req_1;
      type_cast_3327_inst_ack_1<= rack(0);
      type_cast_3327_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3327_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3326_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1518_3328,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3337_inst
    process(add1519_3334) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1519_3334(31 downto 0);
      type_cast_3337_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3339_inst
    process(conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv92_517(31 downto 0);
      type_cast_3339_wire <= tmp_var; -- 
    end process;
    type_cast_3366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3366_inst_req_0;
      type_cast_3366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3366_inst_req_1;
      type_cast_3366_inst_ack_1<= rack(0);
      type_cast_3366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3365_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1533_3367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3375_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3375_inst_req_0;
      type_cast_3375_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3375_inst_req_1;
      type_cast_3375_inst_ack_1<= rack(0);
      type_cast_3375_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3375_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1541_3372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1546_3376,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3392_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3392_inst_req_0;
      type_cast_3392_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3392_inst_req_1;
      type_cast_3392_inst_ack_1<= rack(0);
      type_cast_3392_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3392_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3391_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1549_3393,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3412_inst_req_0;
      type_cast_3412_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3412_inst_req_1;
      type_cast_3412_inst_ack_1<= rack(0);
      type_cast_3412_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3412_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1527_3354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3412_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3416_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3416_inst_req_0;
      type_cast_3416_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3416_inst_req_1;
      type_cast_3416_inst_ack_1<= rack(0);
      type_cast_3416_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3416_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1546x_xi1355x_x2_3381,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3416_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3418_inst_req_0;
      type_cast_3418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3418_inst_req_1;
      type_cast_3418_inst_ack_1<= rack(0);
      type_cast_3418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1355x_x2_3071,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3418_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3422_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3422_inst_req_0;
      type_cast_3422_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3422_inst_req_1;
      type_cast_3422_inst_ack_1<= rack(0);
      type_cast_3422_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3422_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1406x_x2_3388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3422_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3424_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3424_inst_req_0;
      type_cast_3424_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3424_inst_req_1;
      type_cast_3424_inst_ack_1<= rack(0);
      type_cast_3424_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3424_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1406x_x1_3077,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3424_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3445_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3445_inst_req_0;
      type_cast_3445_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3445_inst_req_1;
      type_cast_3445_inst_ack_1<= rack(0);
      type_cast_3445_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3445_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1584_3442,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1635_3446,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_344_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_344_inst_req_0;
      type_cast_344_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_344_inst_req_1;
      type_cast_344_inst_ack_1<= rack(0);
      type_cast_344_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_344_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_495,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_344_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3481_inst_req_0;
      type_cast_3481_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3481_inst_req_1;
      type_cast_3481_inst_ack_1<= rack(0);
      type_cast_3481_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3481_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => k1568x_x0x_xph_3815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3481_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3485_inst_req_0;
      type_cast_3485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3485_inst_req_1;
      type_cast_3485_inst_ack_1<= rack(0);
      type_cast_3485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div1580_3439,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3485_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3487_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3487_inst_req_0;
      type_cast_3487_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3487_inst_req_1;
      type_cast_3487_inst_ack_1<= rack(0);
      type_cast_3487_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3487_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1576x_x1x_xph_3822,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3487_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3491_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3491_inst_req_0;
      type_cast_3491_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3491_inst_req_1;
      type_cast_3491_inst_ack_1<= rack(0);
      type_cast_3491_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3491_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div260_998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3491_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3493_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3493_inst_req_0;
      type_cast_3493_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3493_inst_req_1;
      type_cast_3493_inst_ack_1<= rack(0);
      type_cast_3493_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3493_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1627x_x0x_xph_3828,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3493_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3498_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3498_inst_req_0;
      type_cast_3498_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3498_inst_req_1;
      type_cast_3498_inst_ack_1<= rack(0);
      type_cast_3498_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3498_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3497_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1633_3499,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3502_inst
    process(conv1633_3499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1633_3499(31 downto 0);
      type_cast_3502_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3504_inst
    process(conv1635_3446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1635_3446(31 downto 0);
      type_cast_3504_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3515_inst
    process(conv1633_3499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1633_3499(31 downto 0);
      type_cast_3515_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3517_inst
    process(add1645_3467) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1645_3467(31 downto 0);
      type_cast_3517_wire <= tmp_var; -- 
    end process;
    type_cast_3535_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3535_inst_req_0;
      type_cast_3535_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3535_inst_req_1;
      type_cast_3535_inst_ack_1<= rack(0);
      type_cast_3535_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3535_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3534_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1650_3536,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3539_inst
    process(conv1650_3536) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1650_3536(31 downto 0);
      type_cast_3539_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3541_inst
    process(conv1635_3446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1635_3446(31 downto 0);
      type_cast_3541_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3552_inst
    process(conv1650_3536) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv1650_3536(31 downto 0);
      type_cast_3552_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3554_inst
    process(add1662_3472) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1662_3472(31 downto 0);
      type_cast_3554_wire <= tmp_var; -- 
    end process;
    type_cast_3572_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3572_inst_req_0;
      type_cast_3572_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3572_inst_req_1;
      type_cast_3572_inst_ack_1<= rack(0);
      type_cast_3572_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3572_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3571_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1669_3573,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3577_inst_req_0;
      type_cast_3577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3577_inst_req_1;
      type_cast_3577_inst_ack_1<= rack(0);
      type_cast_3577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3576_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1673_3578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_358_inst_req_0;
      type_cast_358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_358_inst_req_1;
      type_cast_358_inst_ack_1<= rack(0);
      type_cast_358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv21_359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3601_inst
    process(add1681_3598) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1681_3598(31 downto 0);
      type_cast_3601_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3606_inst
    process(ASHR_i32_i32_3605_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3605_wire(31 downto 0);
      shr1683_3607 <= tmp_var; -- 
    end process;
    type_cast_3611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3611_inst_req_0;
      type_cast_3611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3611_inst_req_1;
      type_cast_3611_inst_ack_1<= rack(0);
      type_cast_3611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3610_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1684_3612,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3630_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3630_inst_req_0;
      type_cast_3630_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3630_inst_req_1;
      type_cast_3630_inst_ack_1<= rack(0);
      type_cast_3630_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3630_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3629_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1690_3631,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3684_inst
    process(add1708_3661) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1708_3661(31 downto 0);
      type_cast_3684_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3689_inst
    process(ASHR_i32_i32_3688_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3688_wire(31 downto 0);
      shr1726_3690 <= tmp_var; -- 
    end process;
    type_cast_3694_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3694_inst_req_0;
      type_cast_3694_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3694_inst_req_1;
      type_cast_3694_inst_ack_1<= rack(0);
      type_cast_3694_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3694_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3693_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1727_3695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3709_inst
    process(add1724_3681) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1724_3681(31 downto 0);
      type_cast_3709_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3714_inst
    process(ASHR_i32_i32_3713_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3713_wire(31 downto 0);
      shr1731_3715 <= tmp_var; -- 
    end process;
    type_cast_3719_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3719_inst_req_0;
      type_cast_3719_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3719_inst_req_1;
      type_cast_3719_inst_ack_1<= rack(0);
      type_cast_3719_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3719_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3718_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom1732_3720,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_371_inst_req_0;
      type_cast_371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_371_inst_req_1;
      type_cast_371_inst_ack_1<= rack(0);
      type_cast_371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv25_372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3737_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3737_inst_req_0;
      type_cast_3737_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3737_inst_req_1;
      type_cast_3737_inst_ack_1<= rack(0);
      type_cast_3737_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3737_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3736_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1738_3738,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3747_inst
    process(add1739_3744) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add1739_3744(31 downto 0);
      type_cast_3747_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3749_inst
    process(conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv92_517(31 downto 0);
      type_cast_3749_wire <= tmp_var; -- 
    end process;
    type_cast_3776_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3776_inst_req_0;
      type_cast_3776_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3776_inst_req_1;
      type_cast_3776_inst_ack_1<= rack(0);
      type_cast_3776_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3776_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3775_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1753_3777,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3785_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3785_inst_req_0;
      type_cast_3785_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3785_inst_req_1;
      type_cast_3785_inst_ack_1<= rack(0);
      type_cast_3785_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3785_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp1760_3782,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc1765_3786,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3801_inst_req_0;
      type_cast_3801_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3801_inst_req_1;
      type_cast_3801_inst_ack_1<= rack(0);
      type_cast_3801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3800_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1768_3802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3821_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3821_inst_req_0;
      type_cast_3821_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3821_inst_req_1;
      type_cast_3821_inst_ack_1<= rack(0);
      type_cast_3821_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3821_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add1747_3764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3821_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3825_inst_req_0;
      type_cast_3825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3825_inst_req_1;
      type_cast_3825_inst_ack_1<= rack(0);
      type_cast_3825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i1576x_x2_3482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3825_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3827_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3827_inst_req_0;
      type_cast_3827_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3827_inst_req_1;
      type_cast_3827_inst_ack_1<= rack(0);
      type_cast_3827_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3827_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc1765x_xi1576x_x2_3791,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3827_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3831_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3831_inst_req_0;
      type_cast_3831_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3831_inst_req_1;
      type_cast_3831_inst_ack_1<= rack(0);
      type_cast_3831_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3831_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1627x_x2_3797,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3831_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3833_inst_req_0;
      type_cast_3833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3833_inst_req_1;
      type_cast_3833_inst_ack_1<= rack(0);
      type_cast_3833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => j1627x_x1_3488,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3833_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3840_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3840_inst_req_0;
      type_cast_3840_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3840_inst_req_1;
      type_cast_3840_inst_ack_1<= rack(0);
      type_cast_3840_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3840_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1788_3841,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3844_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3844_inst_req_0;
      type_cast_3844_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3844_inst_req_1;
      type_cast_3844_inst_ack_1<= rack(0);
      type_cast_3844_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3844_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1790_3845,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_389_inst_req_0;
      type_cast_389_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_389_inst_req_1;
      type_cast_389_inst_ack_1<= rack(0);
      type_cast_389_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_386,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_390,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_407_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_407_inst_req_0;
      type_cast_407_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_407_inst_req_1;
      type_cast_407_inst_ack_1<= rack(0);
      type_cast_407_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_407_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call34_404,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_408,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_425_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_425_inst_req_0;
      type_cast_425_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_425_inst_req_1;
      type_cast_425_inst_ack_1<= rack(0);
      type_cast_425_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_425_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call40_422,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_426,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_443_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_443_inst_req_0;
      type_cast_443_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_443_inst_req_1;
      type_cast_443_inst_ack_1<= rack(0);
      type_cast_443_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_443_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_440,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_461_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_461_inst_req_0;
      type_cast_461_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_461_inst_req_1;
      type_cast_461_inst_ack_1<= rack(0);
      type_cast_461_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_461_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call52_458,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv54_462,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_479_inst_req_0;
      type_cast_479_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_479_inst_req_1;
      type_cast_479_inst_ack_1<= rack(0);
      type_cast_479_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_479_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call58_476,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_480,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_516_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_516_inst_req_0;
      type_cast_516_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_516_inst_req_1;
      type_cast_516_inst_ack_1<= rack(0);
      type_cast_516_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_516_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv92_517,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_520_inst_req_0;
      type_cast_520_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_520_inst_req_1;
      type_cast_520_inst_ack_1<= rack(0);
      type_cast_520_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_520_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_524_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_524_inst_req_0;
      type_cast_524_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_524_inst_req_1;
      type_cast_524_inst_ack_1<= rack(0);
      type_cast_524_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_524_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call8_253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_525,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_528_inst_req_0;
      type_cast_528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_528_inst_req_1;
      type_cast_528_inst_ack_1<= rack(0);
      type_cast_528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_537_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_537_inst_req_0;
      type_cast_537_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_537_inst_req_1;
      type_cast_537_inst_ack_1<= rack(0);
      type_cast_537_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_537_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp70_513,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_538,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_541_inst_req_0;
      type_cast_541_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_541_inst_req_1;
      type_cast_541_inst_ack_1<= rack(0);
      type_cast_541_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_541_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call8_253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_542,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_551_inst
    process(sext1848_548) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext1848_548(31 downto 0);
      type_cast_551_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_556_inst
    process(ASHR_i32_i32_555_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_555_wire(31 downto 0);
      conv150_557 <= tmp_var; -- 
    end process;
    type_cast_577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_577_inst_req_0;
      type_cast_577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_577_inst_req_1;
      type_cast_577_inst_ack_1<= rack(0);
      type_cast_577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv239_578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_613_inst
    process(sext_610) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_610(31 downto 0);
      type_cast_613_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_618_inst
    process(ASHR_i32_i32_617_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_617_wire(31 downto 0);
      conv171_619 <= tmp_var; -- 
    end process;
    type_cast_629_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_629_inst_req_0;
      type_cast_629_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_629_inst_req_1;
      type_cast_629_inst_ack_1<= rack(0);
      type_cast_629_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_629_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0x_xph_967,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_629_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_636_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_636_inst_req_0;
      type_cast_636_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_636_inst_req_1;
      type_cast_636_inst_ack_1<= rack(0);
      type_cast_636_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_636_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i68x_x1x_xph_973,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_636_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_643_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_643_inst_req_0;
      type_cast_643_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_643_inst_req_1;
      type_cast_643_inst_ack_1<= rack(0);
      type_cast_643_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_643_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0x_xph_979,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_643_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_648_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_648_inst_req_0;
      type_cast_648_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_648_inst_req_1;
      type_cast_648_inst_ack_1<= rack(0);
      type_cast_648_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_648_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_647_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv108_649,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_652_inst
    process(conv108_649) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv108_649(31 downto 0);
      type_cast_652_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_654_inst
    process(conv110_538) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv110_538(31 downto 0);
      type_cast_654_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_665_inst
    process(conv108_649) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv108_649(31 downto 0);
      type_cast_665_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_667_inst
    process(add119_594) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add119_594(31 downto 0);
      type_cast_667_wire <= tmp_var; -- 
    end process;
    type_cast_685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_685_inst_req_0;
      type_cast_685_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_685_inst_req_1;
      type_cast_685_inst_ack_1<= rack(0);
      type_cast_685_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_685_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_684_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv124_686,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_689_inst
    process(conv124_686) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv124_686(31 downto 0);
      type_cast_689_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_691_inst
    process(conv110_538) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv110_538(31 downto 0);
      type_cast_691_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_702_inst
    process(conv124_686) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv124_686(31 downto 0);
      type_cast_702_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_704_inst
    process(add137_599) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add137_599(31 downto 0);
      type_cast_704_wire <= tmp_var; -- 
    end process;
    type_cast_722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_722_inst_req_0;
      type_cast_722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_722_inst_req_1;
      type_cast_722_inst_ack_1<= rack(0);
      type_cast_722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_721_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv142_723,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_727_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_727_inst_req_0;
      type_cast_727_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_727_inst_req_1;
      type_cast_727_inst_ack_1<= rack(0);
      type_cast_727_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_727_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_726_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv146_728,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_751_inst
    process(add154_748) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add154_748(31 downto 0);
      type_cast_751_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_756_inst
    process(ASHR_i32_i32_755_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_755_wire(31 downto 0);
      shr156_757 <= tmp_var; -- 
    end process;
    type_cast_762_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_762_inst_req_0;
      type_cast_762_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_762_inst_req_1;
      type_cast_762_inst_ack_1<= rack(0);
      type_cast_762_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_762_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_761_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom157_763,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_781_inst_req_0;
      type_cast_781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_781_inst_req_1;
      type_cast_781_inst_ack_1<= rack(0);
      type_cast_781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_781_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_780_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_835_inst
    process(add178_812) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add178_812(31 downto 0);
      type_cast_835_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_840_inst
    process(ASHR_i32_i32_839_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_839_wire(31 downto 0);
      shr196_841 <= tmp_var; -- 
    end process;
    type_cast_845_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_845_inst_req_0;
      type_cast_845_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_845_inst_req_1;
      type_cast_845_inst_ack_1<= rack(0);
      type_cast_845_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_845_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_844_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom197_846,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_860_inst
    process(add194_832) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add194_832(31 downto 0);
      type_cast_860_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_865_inst
    process(ASHR_i32_i32_864_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_864_wire(31 downto 0);
      shr201_866 <= tmp_var; -- 
    end process;
    type_cast_870_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_870_inst_req_0;
      type_cast_870_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_870_inst_req_1;
      type_cast_870_inst_ack_1<= rack(0);
      type_cast_870_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_870_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_869_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom202_871,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_888_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_888_inst_req_0;
      type_cast_888_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_888_inst_req_1;
      type_cast_888_inst_ack_1<= rack(0);
      type_cast_888_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_888_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_887_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_889,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_898_inst
    process(add207_895) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add207_895(31 downto 0);
      type_cast_898_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_900_inst
    process(conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv92_517(31 downto 0);
      type_cast_900_wire <= tmp_var; -- 
    end process;
    type_cast_927_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_927_inst_req_0;
      type_cast_927_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_927_inst_req_1;
      type_cast_927_inst_ack_1<= rack(0);
      type_cast_927_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_927_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_926_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv221_928,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_936_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_936_inst_req_0;
      type_cast_936_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_936_inst_req_1;
      type_cast_936_inst_ack_1<= rack(0);
      type_cast_936_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_936_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp229_933,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc234_937,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_953_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_953_inst_req_0;
      type_cast_953_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_953_inst_req_1;
      type_cast_953_inst_ack_1<= rack(0);
      type_cast_953_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_953_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_952_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv237_954,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_970_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_970_inst_req_0;
      type_cast_970_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_970_inst_req_1;
      type_cast_970_inst_ack_1<= rack(0);
      type_cast_970_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_970_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_622,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_970_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_972_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_972_inst_req_0;
      type_cast_972_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_972_inst_req_1;
      type_cast_972_inst_ack_1<= rack(0);
      type_cast_972_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_972_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_949,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_972_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_976_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_976_inst_req_0;
      type_cast_976_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_976_inst_req_1;
      type_cast_976_inst_ack_1<= rack(0);
      type_cast_976_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_976_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => i68x_x2_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_976_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_978_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_978_inst_req_0;
      type_cast_978_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_978_inst_req_1;
      type_cast_978_inst_ack_1<= rack(0);
      type_cast_978_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_978_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc234x_xi68x_x2_942,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_978_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_982_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_982_inst_req_0;
      type_cast_982_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_982_inst_req_1;
      type_cast_982_inst_ack_1<= rack(0);
      type_cast_982_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_982_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add215_915,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_982_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_991_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_991_inst_req_0;
      type_cast_991_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_991_inst_req_1;
      type_cast_991_inst_ack_1<= rack(0);
      type_cast_991_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_991_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv259_992,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_pad_1000_gather_scatter
    process(LOAD_pad_1000_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_1000_data_0;
      ov(7 downto 0) := iv;
      tmp266_1001 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_1408_gather_scatter
    process(LOAD_pad_1408_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_1408_data_0;
      ov(7 downto 0) := iv;
      tmp482_1409 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_1813_gather_scatter
    process(LOAD_pad_1813_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_1813_data_0;
      ov(7 downto 0) := iv;
      tmp704_1814 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_2216_gather_scatter
    process(LOAD_pad_2216_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_2216_data_0;
      ov(7 downto 0) := iv;
      tmp920_2217 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_2627_gather_scatter
    process(LOAD_pad_2627_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_2627_data_0;
      ov(7 downto 0) := iv;
      tmp1144_2628 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_3030_gather_scatter
    process(LOAD_pad_3030_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_3030_data_0;
      ov(7 downto 0) := iv;
      tmp1363_3031 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_3441_gather_scatter
    process(LOAD_pad_3441_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_3441_data_0;
      ov(7 downto 0) := iv;
      tmp1584_3442 <= ov(7 downto 0);
      --
    end process;
    -- equivalence LOAD_pad_512_gather_scatter
    process(LOAD_pad_512_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_pad_512_data_0;
      ov(7 downto 0) := iv;
      tmp70_513 <= ov(7 downto 0);
      --
    end process;
    -- equivalence STORE_pad_242_gather_scatter
    process(call5_241) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call5_241;
      ov(7 downto 0) := iv;
      STORE_pad_242_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1177_index_1_rename
    process(R_idxprom367_1176_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom367_1176_resized;
      ov(13 downto 0) := iv;
      R_idxprom367_1176_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1177_index_1_resize
    process(idxprom367_1172) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom367_1172;
      ov := iv(13 downto 0);
      R_idxprom367_1176_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1177_root_address_inst
    process(array_obj_ref_1177_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1177_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1177_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1260_index_1_rename
    process(R_idxprom410_1259_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom410_1259_resized;
      ov(13 downto 0) := iv;
      R_idxprom410_1259_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1260_index_1_resize
    process(idxprom410_1255) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom410_1255;
      ov := iv(13 downto 0);
      R_idxprom410_1259_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1260_root_address_inst
    process(array_obj_ref_1260_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1260_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1260_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1285_index_1_rename
    process(R_idxprom415_1284_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom415_1284_resized;
      ov(13 downto 0) := iv;
      R_idxprom415_1284_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1285_index_1_resize
    process(idxprom415_1280) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom415_1280;
      ov := iv(13 downto 0);
      R_idxprom415_1284_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1285_root_address_inst
    process(array_obj_ref_1285_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1285_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1285_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1591_index_1_rename
    process(R_idxprom584_1590_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom584_1590_resized;
      ov(13 downto 0) := iv;
      R_idxprom584_1590_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1591_index_1_resize
    process(idxprom584_1586) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom584_1586;
      ov := iv(13 downto 0);
      R_idxprom584_1590_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1591_root_address_inst
    process(array_obj_ref_1591_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1591_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1591_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1674_index_1_rename
    process(R_idxprom627_1673_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom627_1673_resized;
      ov(13 downto 0) := iv;
      R_idxprom627_1673_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1674_index_1_resize
    process(idxprom627_1669) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom627_1669;
      ov := iv(13 downto 0);
      R_idxprom627_1673_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1674_root_address_inst
    process(array_obj_ref_1674_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1674_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1674_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1699_index_1_rename
    process(R_idxprom632_1698_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom632_1698_resized;
      ov(13 downto 0) := iv;
      R_idxprom632_1698_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1699_index_1_resize
    process(idxprom632_1694) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom632_1694;
      ov := iv(13 downto 0);
      R_idxprom632_1698_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1699_root_address_inst
    process(array_obj_ref_1699_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1699_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1699_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1989_index_1_rename
    process(R_idxprom805_1988_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom805_1988_resized;
      ov(13 downto 0) := iv;
      R_idxprom805_1988_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1989_index_1_resize
    process(idxprom805_1984) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom805_1984;
      ov := iv(13 downto 0);
      R_idxprom805_1988_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1989_root_address_inst
    process(array_obj_ref_1989_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1989_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1989_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2072_index_1_rename
    process(R_idxprom848_2071_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom848_2071_resized;
      ov(13 downto 0) := iv;
      R_idxprom848_2071_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2072_index_1_resize
    process(idxprom848_2067) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom848_2067;
      ov := iv(13 downto 0);
      R_idxprom848_2071_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2072_root_address_inst
    process(array_obj_ref_2072_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2072_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2072_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2097_index_1_rename
    process(R_idxprom853_2096_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom853_2096_resized;
      ov(13 downto 0) := iv;
      R_idxprom853_2096_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2097_index_1_resize
    process(idxprom853_2092) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom853_2092;
      ov := iv(13 downto 0);
      R_idxprom853_2096_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2097_root_address_inst
    process(array_obj_ref_2097_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2097_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2097_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2405_index_1_rename
    process(R_idxprom1023_2404_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1023_2404_resized;
      ov(13 downto 0) := iv;
      R_idxprom1023_2404_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2405_index_1_resize
    process(idxprom1023_2400) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1023_2400;
      ov := iv(13 downto 0);
      R_idxprom1023_2404_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2405_root_address_inst
    process(array_obj_ref_2405_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2405_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2405_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2488_index_1_rename
    process(R_idxprom1066_2487_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1066_2487_resized;
      ov(13 downto 0) := iv;
      R_idxprom1066_2487_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2488_index_1_resize
    process(idxprom1066_2483) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1066_2483;
      ov := iv(13 downto 0);
      R_idxprom1066_2487_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2488_root_address_inst
    process(array_obj_ref_2488_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2488_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2488_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2513_index_1_rename
    process(R_idxprom1071_2512_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1071_2512_resized;
      ov(13 downto 0) := iv;
      R_idxprom1071_2512_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2513_index_1_resize
    process(idxprom1071_2508) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1071_2508;
      ov := iv(13 downto 0);
      R_idxprom1071_2512_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2513_root_address_inst
    process(array_obj_ref_2513_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2513_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2513_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2803_index_1_rename
    process(R_idxprom1246_2802_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1246_2802_resized;
      ov(13 downto 0) := iv;
      R_idxprom1246_2802_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2803_index_1_resize
    process(idxprom1246_2798) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1246_2798;
      ov := iv(13 downto 0);
      R_idxprom1246_2802_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2803_root_address_inst
    process(array_obj_ref_2803_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2803_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2803_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2886_index_1_rename
    process(R_idxprom1289_2885_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1289_2885_resized;
      ov(13 downto 0) := iv;
      R_idxprom1289_2885_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2886_index_1_resize
    process(idxprom1289_2881) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1289_2881;
      ov := iv(13 downto 0);
      R_idxprom1289_2885_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2886_root_address_inst
    process(array_obj_ref_2886_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2886_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2886_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2911_index_1_rename
    process(R_idxprom1294_2910_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1294_2910_resized;
      ov(13 downto 0) := iv;
      R_idxprom1294_2910_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2911_index_1_resize
    process(idxprom1294_2906) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1294_2906;
      ov := iv(13 downto 0);
      R_idxprom1294_2910_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2911_root_address_inst
    process(array_obj_ref_2911_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2911_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2911_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3207_index_1_rename
    process(R_idxprom1464_3206_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1464_3206_resized;
      ov(13 downto 0) := iv;
      R_idxprom1464_3206_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3207_index_1_resize
    process(idxprom1464_3202) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1464_3202;
      ov := iv(13 downto 0);
      R_idxprom1464_3206_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3207_root_address_inst
    process(array_obj_ref_3207_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3207_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3207_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3290_index_1_rename
    process(R_idxprom1507_3289_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1507_3289_resized;
      ov(13 downto 0) := iv;
      R_idxprom1507_3289_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3290_index_1_resize
    process(idxprom1507_3285) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1507_3285;
      ov := iv(13 downto 0);
      R_idxprom1507_3289_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3290_root_address_inst
    process(array_obj_ref_3290_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3290_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3290_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3315_index_1_rename
    process(R_idxprom1512_3314_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1512_3314_resized;
      ov(13 downto 0) := iv;
      R_idxprom1512_3314_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3315_index_1_resize
    process(idxprom1512_3310) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1512_3310;
      ov := iv(13 downto 0);
      R_idxprom1512_3314_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3315_root_address_inst
    process(array_obj_ref_3315_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3315_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3315_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_350_index_1_rename
    process(R_indvar_349_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_349_resized;
      ov(13 downto 0) := iv;
      R_indvar_349_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_350_index_1_resize
    process(indvar_338) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_338;
      ov := iv(13 downto 0);
      R_indvar_349_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_350_root_address_inst
    process(array_obj_ref_350_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_350_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_350_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3617_index_1_rename
    process(R_idxprom1684_3616_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1684_3616_resized;
      ov(13 downto 0) := iv;
      R_idxprom1684_3616_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3617_index_1_resize
    process(idxprom1684_3612) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1684_3612;
      ov := iv(13 downto 0);
      R_idxprom1684_3616_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3617_root_address_inst
    process(array_obj_ref_3617_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3617_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3617_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3700_index_1_rename
    process(R_idxprom1727_3699_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1727_3699_resized;
      ov(13 downto 0) := iv;
      R_idxprom1727_3699_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3700_index_1_resize
    process(idxprom1727_3695) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1727_3695;
      ov := iv(13 downto 0);
      R_idxprom1727_3699_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3700_root_address_inst
    process(array_obj_ref_3700_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3700_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3700_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3725_index_1_rename
    process(R_idxprom1732_3724_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom1732_3724_resized;
      ov(13 downto 0) := iv;
      R_idxprom1732_3724_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3725_index_1_resize
    process(idxprom1732_3720) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom1732_3720;
      ov := iv(13 downto 0);
      R_idxprom1732_3724_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3725_root_address_inst
    process(array_obj_ref_3725_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3725_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3725_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_768_index_1_rename
    process(R_idxprom157_767_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom157_767_resized;
      ov(13 downto 0) := iv;
      R_idxprom157_767_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_768_index_1_resize
    process(idxprom157_763) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom157_763;
      ov := iv(13 downto 0);
      R_idxprom157_767_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_768_root_address_inst
    process(array_obj_ref_768_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_768_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_768_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_851_index_1_rename
    process(R_idxprom197_850_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom197_850_resized;
      ov(13 downto 0) := iv;
      R_idxprom197_850_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_851_index_1_resize
    process(idxprom197_846) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom197_846;
      ov := iv(13 downto 0);
      R_idxprom197_850_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_851_root_address_inst
    process(array_obj_ref_851_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_851_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_851_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_index_1_rename
    process(R_idxprom202_875_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom202_875_resized;
      ov(13 downto 0) := iv;
      R_idxprom202_875_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_index_1_resize
    process(idxprom202_871) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom202_871;
      ov := iv(13 downto 0);
      R_idxprom202_875_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_root_address_inst
    process(array_obj_ref_876_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_876_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_876_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1181_addr_0
    process(ptr_deref_1181_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1181_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1181_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1181_base_resize
    process(arrayidx368_1179) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx368_1179;
      ov := iv(13 downto 0);
      ptr_deref_1181_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1181_gather_scatter
    process(type_cast_1183_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1183_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1181_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1181_root_address_inst
    process(ptr_deref_1181_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1181_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1181_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1265_addr_0
    process(ptr_deref_1265_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1265_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1265_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1265_base_resize
    process(arrayidx411_1262) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx411_1262;
      ov := iv(13 downto 0);
      ptr_deref_1265_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1265_gather_scatter
    process(ptr_deref_1265_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1265_data_0;
      ov(63 downto 0) := iv;
      tmp412_1266 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1265_root_address_inst
    process(ptr_deref_1265_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1265_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1265_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1289_addr_0
    process(ptr_deref_1289_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1289_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1289_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1289_base_resize
    process(arrayidx416_1287) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx416_1287;
      ov := iv(13 downto 0);
      ptr_deref_1289_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1289_gather_scatter
    process(tmp412_1266) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp412_1266;
      ov(63 downto 0) := iv;
      ptr_deref_1289_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1289_root_address_inst
    process(ptr_deref_1289_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1289_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1289_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1595_addr_0
    process(ptr_deref_1595_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1595_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1595_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1595_base_resize
    process(arrayidx585_1593) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx585_1593;
      ov := iv(13 downto 0);
      ptr_deref_1595_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1595_gather_scatter
    process(type_cast_1597_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1597_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1595_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1595_root_address_inst
    process(ptr_deref_1595_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1595_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1595_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1679_addr_0
    process(ptr_deref_1679_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1679_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1679_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1679_base_resize
    process(arrayidx628_1676) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx628_1676;
      ov := iv(13 downto 0);
      ptr_deref_1679_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1679_gather_scatter
    process(ptr_deref_1679_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1679_data_0;
      ov(63 downto 0) := iv;
      tmp629_1680 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1679_root_address_inst
    process(ptr_deref_1679_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1679_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1679_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1703_addr_0
    process(ptr_deref_1703_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1703_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1703_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1703_base_resize
    process(arrayidx633_1701) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx633_1701;
      ov := iv(13 downto 0);
      ptr_deref_1703_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1703_gather_scatter
    process(tmp629_1680) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp629_1680;
      ov(63 downto 0) := iv;
      ptr_deref_1703_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1703_root_address_inst
    process(ptr_deref_1703_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1703_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1703_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1993_addr_0
    process(ptr_deref_1993_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1993_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1993_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1993_base_resize
    process(arrayidx806_1991) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx806_1991;
      ov := iv(13 downto 0);
      ptr_deref_1993_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1993_gather_scatter
    process(type_cast_1995_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1995_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1993_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1993_root_address_inst
    process(ptr_deref_1993_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1993_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1993_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2077_addr_0
    process(ptr_deref_2077_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2077_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2077_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2077_base_resize
    process(arrayidx849_2074) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx849_2074;
      ov := iv(13 downto 0);
      ptr_deref_2077_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2077_gather_scatter
    process(ptr_deref_2077_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2077_data_0;
      ov(63 downto 0) := iv;
      tmp850_2078 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2077_root_address_inst
    process(ptr_deref_2077_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2077_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2077_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_addr_0
    process(ptr_deref_2101_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2101_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2101_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_base_resize
    process(arrayidx854_2099) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx854_2099;
      ov := iv(13 downto 0);
      ptr_deref_2101_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_gather_scatter
    process(tmp850_2078) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp850_2078;
      ov(63 downto 0) := iv;
      ptr_deref_2101_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2101_root_address_inst
    process(ptr_deref_2101_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2101_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2101_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2409_addr_0
    process(ptr_deref_2409_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2409_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2409_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2409_base_resize
    process(arrayidx1024_2407) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1024_2407;
      ov := iv(13 downto 0);
      ptr_deref_2409_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2409_gather_scatter
    process(type_cast_2411_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2411_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2409_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2409_root_address_inst
    process(ptr_deref_2409_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2409_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2409_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2493_addr_0
    process(ptr_deref_2493_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2493_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2493_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2493_base_resize
    process(arrayidx1067_2490) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1067_2490;
      ov := iv(13 downto 0);
      ptr_deref_2493_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2493_gather_scatter
    process(ptr_deref_2493_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2493_data_0;
      ov(63 downto 0) := iv;
      tmp1068_2494 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2493_root_address_inst
    process(ptr_deref_2493_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2493_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2493_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2517_addr_0
    process(ptr_deref_2517_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2517_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2517_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2517_base_resize
    process(arrayidx1072_2515) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1072_2515;
      ov := iv(13 downto 0);
      ptr_deref_2517_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2517_gather_scatter
    process(tmp1068_2494) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1068_2494;
      ov(63 downto 0) := iv;
      ptr_deref_2517_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2517_root_address_inst
    process(ptr_deref_2517_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2517_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2517_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2807_addr_0
    process(ptr_deref_2807_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2807_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2807_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2807_base_resize
    process(arrayidx1247_2805) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1247_2805;
      ov := iv(13 downto 0);
      ptr_deref_2807_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2807_gather_scatter
    process(type_cast_2809_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2809_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2807_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2807_root_address_inst
    process(ptr_deref_2807_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2807_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2807_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2891_addr_0
    process(ptr_deref_2891_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2891_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2891_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2891_base_resize
    process(arrayidx1290_2888) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1290_2888;
      ov := iv(13 downto 0);
      ptr_deref_2891_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2891_gather_scatter
    process(ptr_deref_2891_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2891_data_0;
      ov(63 downto 0) := iv;
      tmp1291_2892 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2891_root_address_inst
    process(ptr_deref_2891_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2891_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2891_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2915_addr_0
    process(ptr_deref_2915_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2915_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2915_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2915_base_resize
    process(arrayidx1295_2913) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1295_2913;
      ov := iv(13 downto 0);
      ptr_deref_2915_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2915_gather_scatter
    process(tmp1291_2892) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1291_2892;
      ov(63 downto 0) := iv;
      ptr_deref_2915_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2915_root_address_inst
    process(ptr_deref_2915_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2915_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2915_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3211_addr_0
    process(ptr_deref_3211_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3211_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3211_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3211_base_resize
    process(arrayidx1465_3209) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1465_3209;
      ov := iv(13 downto 0);
      ptr_deref_3211_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3211_gather_scatter
    process(type_cast_3213_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3213_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3211_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3211_root_address_inst
    process(ptr_deref_3211_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3211_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3211_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3295_addr_0
    process(ptr_deref_3295_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3295_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3295_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3295_base_resize
    process(arrayidx1508_3292) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1508_3292;
      ov := iv(13 downto 0);
      ptr_deref_3295_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3295_gather_scatter
    process(ptr_deref_3295_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3295_data_0;
      ov(63 downto 0) := iv;
      tmp1509_3296 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3295_root_address_inst
    process(ptr_deref_3295_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3295_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3295_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3319_addr_0
    process(ptr_deref_3319_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3319_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3319_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3319_base_resize
    process(arrayidx1513_3317) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1513_3317;
      ov := iv(13 downto 0);
      ptr_deref_3319_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3319_gather_scatter
    process(tmp1509_3296) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1509_3296;
      ov(63 downto 0) := iv;
      ptr_deref_3319_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3319_root_address_inst
    process(ptr_deref_3319_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3319_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3319_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3621_addr_0
    process(ptr_deref_3621_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3621_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3621_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3621_base_resize
    process(arrayidx1685_3619) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1685_3619;
      ov := iv(13 downto 0);
      ptr_deref_3621_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3621_gather_scatter
    process(type_cast_3623_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3623_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_3621_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3621_root_address_inst
    process(ptr_deref_3621_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3621_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3621_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3705_addr_0
    process(ptr_deref_3705_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3705_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3705_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3705_base_resize
    process(arrayidx1728_3702) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1728_3702;
      ov := iv(13 downto 0);
      ptr_deref_3705_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3705_gather_scatter
    process(ptr_deref_3705_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3705_data_0;
      ov(63 downto 0) := iv;
      tmp1729_3706 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3705_root_address_inst
    process(ptr_deref_3705_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3705_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3705_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3729_addr_0
    process(ptr_deref_3729_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3729_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3729_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3729_base_resize
    process(arrayidx1733_3727) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx1733_3727;
      ov := iv(13 downto 0);
      ptr_deref_3729_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3729_gather_scatter
    process(tmp1729_3706) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp1729_3706;
      ov(63 downto 0) := iv;
      ptr_deref_3729_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3729_root_address_inst
    process(ptr_deref_3729_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3729_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3729_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_487_addr_0
    process(ptr_deref_487_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_487_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_487_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_487_base_resize
    process(arrayidx_352) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_352;
      ov := iv(13 downto 0);
      ptr_deref_487_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_487_gather_scatter
    process(add61_485) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add61_485;
      ov(63 downto 0) := iv;
      ptr_deref_487_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_487_root_address_inst
    process(ptr_deref_487_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_487_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_487_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_772_addr_0
    process(ptr_deref_772_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_772_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_772_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_772_base_resize
    process(arrayidx158_770) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx158_770;
      ov := iv(13 downto 0);
      ptr_deref_772_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_772_gather_scatter
    process(type_cast_774_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_774_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_772_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_772_root_address_inst
    process(ptr_deref_772_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_772_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_772_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_856_addr_0
    process(ptr_deref_856_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_856_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_856_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_856_base_resize
    process(arrayidx198_853) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx198_853;
      ov := iv(13 downto 0);
      ptr_deref_856_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_856_gather_scatter
    process(ptr_deref_856_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_856_data_0;
      ov(63 downto 0) := iv;
      tmp199_857 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_856_root_address_inst
    process(ptr_deref_856_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_856_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_856_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_addr_0
    process(ptr_deref_880_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_880_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_880_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_base_resize
    process(arrayidx203_878) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx203_878;
      ov := iv(13 downto 0);
      ptr_deref_880_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_gather_scatter
    process(tmp199_857) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp199_857;
      ov(63 downto 0) := iv;
      ptr_deref_880_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_880_root_address_inst
    process(ptr_deref_880_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_880_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_880_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1085_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1850_1084;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1085_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1085_branch_req_0,
          ack0 => if_stmt_1085_branch_ack_0,
          ack1 => if_stmt_1085_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1122_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1851_1121;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1122_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1122_branch_req_0,
          ack0 => if_stmt_1122_branch_ack_0,
          ack1 => if_stmt_1122_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1312_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp425_1311;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1312_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1312_branch_req_0,
          ack0 => if_stmt_1312_branch_ack_0,
          ack1 => if_stmt_1312_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1368_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp459_1367;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1368_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1368_branch_req_0,
          ack0 => if_stmt_1368_branch_ack_0,
          ack1 => if_stmt_1368_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1499_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1852_1498;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1499_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1499_branch_req_0,
          ack0 => if_stmt_1499_branch_ack_0,
          ack1 => if_stmt_1499_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1536_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1853_1535;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1536_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1536_branch_req_0,
          ack0 => if_stmt_1536_branch_ack_0,
          ack1 => if_stmt_1536_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1726_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp642_1725;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1726_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1726_branch_req_0,
          ack0 => if_stmt_1726_branch_ack_0,
          ack1 => if_stmt_1726_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1783_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp677_1782;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1783_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1783_branch_req_0,
          ack0 => if_stmt_1783_branch_ack_0,
          ack1 => if_stmt_1783_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1897_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1854_1896;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1897_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1897_branch_req_0,
          ack0 => if_stmt_1897_branch_ack_0,
          ack1 => if_stmt_1897_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1934_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1855_1933;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1934_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1934_branch_req_0,
          ack0 => if_stmt_1934_branch_ack_0,
          ack1 => if_stmt_1934_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2124_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp863_2123;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2124_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2124_branch_req_0,
          ack0 => if_stmt_2124_branch_ack_0,
          ack1 => if_stmt_2124_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2180_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp897_2179;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2180_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2180_branch_req_0,
          ack0 => if_stmt_2180_branch_ack_0,
          ack1 => if_stmt_2180_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2313_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1856_2312;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2313_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2313_branch_req_0,
          ack0 => if_stmt_2313_branch_ack_0,
          ack1 => if_stmt_2313_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2350_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1857_2349;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2350_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2350_branch_req_0,
          ack0 => if_stmt_2350_branch_ack_0,
          ack1 => if_stmt_2350_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2540_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1081_2539;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2540_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2540_branch_req_0,
          ack0 => if_stmt_2540_branch_ack_0,
          ack1 => if_stmt_2540_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2597_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1117_2596;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2597_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2597_branch_req_0,
          ack0 => if_stmt_2597_branch_ack_0,
          ack1 => if_stmt_2597_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2711_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1858_2710;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2711_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2711_branch_req_0,
          ack0 => if_stmt_2711_branch_ack_0,
          ack1 => if_stmt_2711_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2748_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1859_2747;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2748_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2748_branch_req_0,
          ack0 => if_stmt_2748_branch_ack_0,
          ack1 => if_stmt_2748_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_288_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1840_287;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_288_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_288_branch_req_0,
          ack0 => if_stmt_288_branch_ack_0,
          ack1 => if_stmt_288_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2938_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1304_2937;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2938_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2938_branch_req_0,
          ack0 => if_stmt_2938_branch_ack_0,
          ack1 => if_stmt_2938_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2994_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1339_2993;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2994_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2994_branch_req_0,
          ack0 => if_stmt_2994_branch_ack_0,
          ack1 => if_stmt_2994_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3115_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1860_3114;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3115_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3115_branch_req_0,
          ack0 => if_stmt_3115_branch_ack_0,
          ack1 => if_stmt_3115_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3152_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1861_3151;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3152_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3152_branch_req_0,
          ack0 => if_stmt_3152_branch_ack_0,
          ack1 => if_stmt_3152_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3342_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1522_3341;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3342_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3342_branch_req_0,
          ack0 => if_stmt_3342_branch_ack_0,
          ack1 => if_stmt_3342_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3399_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1556_3398;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3399_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3399_branch_req_0,
          ack0 => if_stmt_3399_branch_ack_0,
          ack1 => if_stmt_3399_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3525_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1862_3524;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3525_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3525_branch_req_0,
          ack0 => if_stmt_3525_branch_ack_0,
          ack1 => if_stmt_3525_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3562_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1863_3561;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3562_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3562_branch_req_0,
          ack0 => if_stmt_3562_branch_ack_0,
          ack1 => if_stmt_3562_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3752_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1742_3751;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3752_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3752_branch_req_0,
          ack0 => if_stmt_3752_branch_ack_0,
          ack1 => if_stmt_3752_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3808_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp1775_3807;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3808_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3808_branch_req_0,
          ack0 => if_stmt_3808_branch_ack_0,
          ack1 => if_stmt_3808_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_501_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond8_500;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_501_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_501_branch_req_0,
          ack0 => if_stmt_501_branch_ack_0,
          ack1 => if_stmt_501_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_675_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond_674;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_675_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_675_branch_req_0,
          ack0 => if_stmt_675_branch_ack_0,
          ack1 => if_stmt_675_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_712_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcond1849_711;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_712_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_712_branch_req_0,
          ack0 => if_stmt_712_branch_ack_0,
          ack1 => if_stmt_712_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_903_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp210_902;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_903_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_903_branch_req_0,
          ack0 => if_stmt_903_branch_ack_0,
          ack1 => if_stmt_903_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_960_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp245_959;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_960_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_960_branch_req_0,
          ack0 => if_stmt_960_branch_ack_0,
          ack1 => if_stmt_960_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1323_inst
    process(k255x_x1_1047) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k255x_x1_1047, type_cast_1322_wire_constant, tmp_var);
      add430_1324 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1331_inst
    process(j309x_x1_1034) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j309x_x1_1034, type_cast_1330_wire_constant, tmp_var);
      inc434_1332 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1350_inst
    process(inc448_1346, i263x_x2_1040) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc448_1346, i263x_x2_1040, tmp_var);
      inc448x_xi263x_x2_1351 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1737_inst
    process(k471x_x1_1448) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k471x_x1_1448, type_cast_1736_wire_constant, tmp_var);
      add647_1738 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1745_inst
    process(j525x_x1_1461) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j525x_x1_1461, type_cast_1744_wire_constant, tmp_var);
      inc651_1746 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1764_inst
    process(inc666_1760, i475x_x2_1455) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc666_1760, i475x_x2_1455, tmp_var);
      inc666x_xi475x_x2_1765 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2135_inst
    process(k689x_x1_1847) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k689x_x1_1847, type_cast_2134_wire_constant, tmp_var);
      add868_2136 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2143_inst
    process(j747x_x1_1860) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j747x_x1_1860, type_cast_2142_wire_constant, tmp_var);
      inc872_2144 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2162_inst
    process(inc886_2158, i697x_x2_1854) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc886_2158, i697x_x2_1854, tmp_var);
      inc886x_xi697x_x2_2163 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2551_inst
    process(k909x_x1_2262) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k909x_x1_2262, type_cast_2550_wire_constant, tmp_var);
      add1086_2552 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2559_inst
    process(j963x_x1_2275) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j963x_x1_2275, type_cast_2558_wire_constant, tmp_var);
      inc1090_2560 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2578_inst
    process(inc1105_2574, i913x_x2_2269) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1105_2574, i913x_x2_2269, tmp_var);
      inc1105x_xi913x_x2_2579 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2949_inst
    process(k1129x_x1_2661) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1129x_x1_2661, type_cast_2948_wire_constant, tmp_var);
      add1309_2950 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2957_inst
    process(j1187x_x1_2674) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1187x_x1_2674, type_cast_2956_wire_constant, tmp_var);
      inc1313_2958 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2976_inst
    process(inc1327_2972, i1137x_x2_2668) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1327_2972, i1137x_x2_2668, tmp_var);
      inc1327x_xi1137x_x2_2977 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3353_inst
    process(k1351x_x1_3064) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1351x_x1_3064, type_cast_3352_wire_constant, tmp_var);
      add1527_3354 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3361_inst
    process(j1406x_x1_3077) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1406x_x1_3077, type_cast_3360_wire_constant, tmp_var);
      inc1531_3362 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3380_inst
    process(inc1546_3376, i1355x_x2_3071) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1546_3376, i1355x_x2_3071, tmp_var);
      inc1546x_xi1355x_x2_3381 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3763_inst
    process(k1568x_x1_3475) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(k1568x_x1_3475, type_cast_3762_wire_constant, tmp_var);
      add1747_3764 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3771_inst
    process(j1627x_x1_3488) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(j1627x_x1_3488, type_cast_3770_wire_constant, tmp_var);
      inc1751_3772 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3790_inst
    process(inc1765_3786, i1576x_x2_3482) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc1765_3786, i1576x_x2_3482, tmp_var);
      inc1765x_xi1576x_x2_3791 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_914_inst
    process(kx_x1_637) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_637, type_cast_913_wire_constant, tmp_var);
      add215_915 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_922_inst
    process(jx_x1_622) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_622, type_cast_921_wire_constant, tmp_var);
      inc219_923 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_941_inst
    process(inc234_937, i68x_x2_630) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc234_937, i68x_x2_630, tmp_var);
      inc234x_xi68x_x2_942 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1015_inst
    process(shl441_1011, conv94_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl441_1011, conv94_521, tmp_var);
      add442_1016 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1020_inst
    process(shl441_1011, div240_584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl441_1011, div240_584, tmp_var);
      add458_1021 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1025_inst
    process(conv317_1005, div240_584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv317_1005, div240_584, tmp_var);
      add328_1026 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1030_inst
    process(conv317_1005, conv94_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv317_1005, conv94_521, tmp_var);
      add345_1031 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1152_inst
    process(mul363_1148, mul357_1143) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul363_1148, mul357_1143, tmp_var);
      add358_1153 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1157_inst
    process(add358_1153, conv352_1133) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add358_1153, conv352_1133, tmp_var);
      add364_1158 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1215_inst
    process(conv373_1191, mul381_1201) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv373_1191, mul381_1201, tmp_var);
      add382_1216 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1220_inst
    process(add382_1216, mul390_1211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add382_1216, mul390_1211, tmp_var);
      add391_1221 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1235_inst
    process(mul406_1231, mul400_1226) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul406_1231, mul400_1226, tmp_var);
      add401_1236 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1240_inst
    process(add401_1236, conv373_1191) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add401_1236, conv373_1191, tmp_var);
      add407_1241 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1303_inst
    process(conv421_1298) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv421_1298, type_cast_1302_wire_constant, tmp_var);
      add422_1304 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1423_inst
    process(shl659_1419, div224_563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl659_1419, div224_563, tmp_var);
      add660_1424 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1434_inst
    process(shl659_1419, div672_1430) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl659_1419, div672_1430, tmp_var);
      add676_1435 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1439_inst
    process(conv533_1413, div672_1430) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv533_1413, div672_1430, tmp_var);
      add544_1440 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1444_inst
    process(conv533_1413, div224_563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv533_1413, div224_563, tmp_var);
      add562_1445 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1566_inst
    process(mul580_1562, conv569_1547) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul580_1562, conv569_1547, tmp_var);
      add575_1567 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1571_inst
    process(add575_1567, mul574_1557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add575_1567, mul574_1557, tmp_var);
      add581_1572 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1629_inst
    process(mul607_1625, conv590_1605) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul607_1625, conv590_1605, tmp_var);
      add599_1630 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1634_inst
    process(add599_1630, mul598_1615) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add599_1630, mul598_1615, tmp_var);
      add608_1635 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1649_inst
    process(mul623_1645, conv590_1605) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul623_1645, conv590_1605, tmp_var);
      add618_1650 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1654_inst
    process(add618_1650, mul617_1640) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add618_1650, mul617_1640, tmp_var);
      add624_1655 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1717_inst
    process(conv638_1712) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv638_1712, type_cast_1716_wire_constant, tmp_var);
      add639_1718 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1828_inst
    process(shl879_1824, conv94_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl879_1824, conv94_521, tmp_var);
      add880_1829 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1833_inst
    process(shl879_1824, div672_1430) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl879_1824, div672_1430, tmp_var);
      add896_1834 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1838_inst
    process(conv755_1818, div672_1430) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv755_1818, div672_1430, tmp_var);
      add766_1839 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1843_inst
    process(conv755_1818, conv94_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv755_1818, conv94_521, tmp_var);
      add783_1844 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1964_inst
    process(mul801_1960, conv790_1945) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul801_1960, conv790_1945, tmp_var);
      add796_1965 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1969_inst
    process(add796_1965, mul795_1955) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add796_1965, mul795_1955, tmp_var);
      add802_1970 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2027_inst
    process(mul828_2023, conv811_2003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul828_2023, conv811_2003, tmp_var);
      add820_2028 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2032_inst
    process(add820_2028, mul819_2013) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add820_2028, mul819_2013, tmp_var);
      add829_2033 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2047_inst
    process(mul844_2043, conv811_2003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul844_2043, conv811_2003, tmp_var);
      add839_2048 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2052_inst
    process(add839_2048, mul838_2038) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add839_2048, mul838_2038, tmp_var);
      add845_2053 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2115_inst
    process(conv859_2110) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv859_2110, type_cast_2114_wire_constant, tmp_var);
      add860_2116 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2231_inst
    process(shl1098_2227, div224_563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl1098_2227, div224_563, tmp_var);
      add1099_2232 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2248_inst
    process(shl1098_2227, div1112_2244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl1098_2227, div1112_2244, tmp_var);
      add1116_2249 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2253_inst
    process(conv971_2221, div1112_2244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv971_2221, div1112_2244, tmp_var);
      add983_2254 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2258_inst
    process(conv971_2221, div224_563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv971_2221, div224_563, tmp_var);
      add1001_2259 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2380_inst
    process(mul1019_2376, conv1008_2361) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1019_2376, conv1008_2361, tmp_var);
      add1014_2381 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2385_inst
    process(add1014_2381, mul1013_2371) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1014_2381, mul1013_2371, tmp_var);
      add1020_2386 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2443_inst
    process(mul1046_2439, conv1029_2419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1046_2439, conv1029_2419, tmp_var);
      add1038_2444 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2448_inst
    process(add1038_2444, mul1037_2429) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1038_2444, mul1037_2429, tmp_var);
      add1047_2449 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2463_inst
    process(mul1062_2459, conv1029_2419) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1062_2459, conv1029_2419, tmp_var);
      add1057_2464 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2468_inst
    process(add1057_2464, mul1056_2454) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1057_2464, mul1056_2454, tmp_var);
      add1063_2469 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2531_inst
    process(conv1077_2526) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1077_2526, type_cast_2530_wire_constant, tmp_var);
      add1078_2532 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2642_inst
    process(shl1320_2638, conv94_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl1320_2638, conv94_521, tmp_var);
      add1321_2643 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2647_inst
    process(shl1320_2638, div1112_2244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl1320_2638, div1112_2244, tmp_var);
      add1338_2648 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2652_inst
    process(conv1195_2632, div1112_2244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1195_2632, div1112_2244, tmp_var);
      add1207_2653 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2657_inst
    process(conv1195_2632, conv94_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1195_2632, conv94_521, tmp_var);
      add1224_2658 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2778_inst
    process(mul1242_2774, conv1231_2759) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1242_2774, conv1231_2759, tmp_var);
      add1237_2779 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2783_inst
    process(add1237_2779, mul1236_2769) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1237_2779, mul1236_2769, tmp_var);
      add1243_2784 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2841_inst
    process(mul1269_2837, conv1252_2817) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1269_2837, conv1252_2817, tmp_var);
      add1261_2842 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2846_inst
    process(add1261_2842, mul1260_2827) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1261_2842, mul1260_2827, tmp_var);
      add1270_2847 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2861_inst
    process(mul1285_2857, conv1252_2817) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1285_2857, conv1252_2817, tmp_var);
      add1280_2862 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2866_inst
    process(add1280_2862, mul1279_2852) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1280_2862, mul1279_2852, tmp_var);
      add1286_2867 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2929_inst
    process(conv1300_2924) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1300_2924, type_cast_2928_wire_constant, tmp_var);
      add1301_2930 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3045_inst
    process(shl1539_3041, div224_563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl1539_3041, div224_563, tmp_var);
      add1540_3046 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3050_inst
    process(shl1539_3041, conv239_578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl1539_3041, conv239_578, tmp_var);
      add1555_3051 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3055_inst
    process(conv1414_3035, conv239_578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1414_3035, conv239_578, tmp_var);
      add1424_3056 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3060_inst
    process(conv1414_3035, div224_563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1414_3035, div224_563, tmp_var);
      add1442_3061 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3182_inst
    process(mul1460_3178, conv1449_3163) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1460_3178, conv1449_3163, tmp_var);
      add1455_3183 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3187_inst
    process(add1455_3183, mul1454_3173) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1455_3183, mul1454_3173, tmp_var);
      add1461_3188 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3245_inst
    process(mul1487_3241, conv1470_3221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1487_3241, conv1470_3221, tmp_var);
      add1479_3246 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3250_inst
    process(add1479_3246, mul1478_3231) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1479_3246, mul1478_3231, tmp_var);
      add1488_3251 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3265_inst
    process(mul1503_3261, conv1470_3221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1503_3261, conv1470_3221, tmp_var);
      add1498_3266 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3270_inst
    process(add1498_3266, mul1497_3256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1498_3266, mul1497_3256, tmp_var);
      add1504_3271 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3333_inst
    process(conv1518_3328) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1518_3328, type_cast_3332_wire_constant, tmp_var);
      add1519_3334 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3456_inst
    process(shl1758_3452, conv94_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl1758_3452, conv94_521, tmp_var);
      add1759_3457 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3461_inst
    process(shl1758_3452, conv239_578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl1758_3452, conv239_578, tmp_var);
      add1774_3462 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3466_inst
    process(conv1635_3446, conv239_578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1635_3446, conv239_578, tmp_var);
      add1645_3467 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3471_inst
    process(conv1635_3446, conv94_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1635_3446, conv94_521, tmp_var);
      add1662_3472 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3592_inst
    process(mul1680_3588, conv1669_3573) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1680_3588, conv1669_3573, tmp_var);
      add1675_3593 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3597_inst
    process(add1675_3593, mul1674_3583) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1675_3593, mul1674_3583, tmp_var);
      add1681_3598 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3655_inst
    process(mul1707_3651, conv1690_3631) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1707_3651, conv1690_3631, tmp_var);
      add1699_3656 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3660_inst
    process(add1699_3656, mul1698_3641) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1699_3656, mul1698_3641, tmp_var);
      add1708_3661 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3675_inst
    process(mul1723_3671, conv1690_3631) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul1723_3671, conv1690_3631, tmp_var);
      add1718_3676 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3680_inst
    process(add1718_3676, mul1717_3666) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add1718_3676, mul1717_3666, tmp_var);
      add1724_3681 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3743_inst
    process(conv1738_3738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv1738_3738, type_cast_3742_wire_constant, tmp_var);
      add1739_3744 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_573_inst
    process(shl227_569, div224_563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl227_569, div224_563, tmp_var);
      add228_574 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_588_inst
    process(shl227_569, div240_584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl227_569, div240_584, tmp_var);
      add244_589 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_593_inst
    process(conv110_538, div240_584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv110_538, div240_584, tmp_var);
      add119_594 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_598_inst
    process(conv110_538, div224_563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv110_538, div224_563, tmp_var);
      add137_599 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_742_inst
    process(mul153_738, mul147_733) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul153_738, mul147_733, tmp_var);
      add148_743 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_747_inst
    process(add148_743, conv142_723) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add148_743, conv142_723, tmp_var);
      add154_748 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_806_inst
    process(conv161_782, mul168_792) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv161_782, mul168_792, tmp_var);
      add169_807 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_811_inst
    process(add169_807, mul177_802) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add169_807, mul177_802, tmp_var);
      add178_812 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_826_inst
    process(mul193_822, mul187_817) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul193_822, mul187_817, tmp_var);
      add188_827 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_831_inst
    process(add188_827, conv161_782) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add188_827, conv161_782, tmp_var);
      add194_832 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_894_inst
    process(conv206_889) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv206_889, type_cast_893_wire_constant, tmp_var);
      add207_895 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_494_inst
    process(indvar_338) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_338, type_cast_493_wire_constant, tmp_var);
      indvarx_xnext_495 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1083_inst
    process(cmp318x_xnot_1072, cmp329_1079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp318x_xnot_1072, cmp329_1079, tmp_var);
      orx_xcond1850_1084 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1120_inst
    process(cmp336x_xnot_1109, cmp346_1116) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp336x_xnot_1109, cmp346_1116, tmp_var);
      orx_xcond1851_1121 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1497_inst
    process(cmp534x_xnot_1486, cmp545_1493) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp534x_xnot_1486, cmp545_1493, tmp_var);
      orx_xcond1852_1498 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1534_inst
    process(cmp552x_xnot_1523, cmp563_1530) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp552x_xnot_1523, cmp563_1530, tmp_var);
      orx_xcond1853_1535 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1895_inst
    process(cmp756x_xnot_1884, cmp767_1891) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp756x_xnot_1884, cmp767_1891, tmp_var);
      orx_xcond1854_1896 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1932_inst
    process(cmp774x_xnot_1921, cmp784_1928) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp774x_xnot_1921, cmp784_1928, tmp_var);
      orx_xcond1855_1933 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2311_inst
    process(cmp972x_xnot_2300, cmp984_2307) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp972x_xnot_2300, cmp984_2307, tmp_var);
      orx_xcond1856_2312 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2348_inst
    process(cmp991x_xnot_2337, cmp1002_2344) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp991x_xnot_2337, cmp1002_2344, tmp_var);
      orx_xcond1857_2349 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2709_inst
    process(cmp1196x_xnot_2698, cmp1208_2705) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp1196x_xnot_2698, cmp1208_2705, tmp_var);
      orx_xcond1858_2710 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2746_inst
    process(cmp1215x_xnot_2735, cmp1225_2742) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp1215x_xnot_2735, cmp1225_2742, tmp_var);
      orx_xcond1859_2747 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3113_inst
    process(cmp1415x_xnot_3102, cmp1425_3109) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp1415x_xnot_3102, cmp1425_3109, tmp_var);
      orx_xcond1860_3114 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3150_inst
    process(cmp1432x_xnot_3139, cmp1443_3146) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp1432x_xnot_3139, cmp1443_3146, tmp_var);
      orx_xcond1861_3151 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3523_inst
    process(cmp1636x_xnot_3512, cmp1646_3519) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp1636x_xnot_3512, cmp1646_3519, tmp_var);
      orx_xcond1862_3524 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3560_inst
    process(cmp1653x_xnot_3549, cmp1663_3556) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp1653x_xnot_3549, cmp1663_3556, tmp_var);
      orx_xcond1863_3561 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_673_inst
    process(cmp111x_xnot_662, cmp120_669) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp111x_xnot_662, cmp120_669, tmp_var);
      orx_xcond_674 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_710_inst
    process(cmp127x_xnot_699, cmp138_706) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp127x_xnot_699, cmp138_706, tmp_var);
      orx_xcond1849_711 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_280_inst
    process(mul13_275) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul13_275, type_cast_279_wire_constant, tmp_var);
      shr1839x_xmask_281 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1165_inst
    process(type_cast_1161_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1161_wire, type_cast_1164_wire_constant, tmp_var);
      ASHR_i32_i32_1165_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1248_inst
    process(type_cast_1244_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1244_wire, type_cast_1247_wire_constant, tmp_var);
      ASHR_i32_i32_1248_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1273_inst
    process(type_cast_1269_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1269_wire, type_cast_1272_wire_constant, tmp_var);
      ASHR_i32_i32_1273_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1579_inst
    process(type_cast_1575_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1575_wire, type_cast_1578_wire_constant, tmp_var);
      ASHR_i32_i32_1579_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1662_inst
    process(type_cast_1658_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1658_wire, type_cast_1661_wire_constant, tmp_var);
      ASHR_i32_i32_1662_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1687_inst
    process(type_cast_1683_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1683_wire, type_cast_1686_wire_constant, tmp_var);
      ASHR_i32_i32_1687_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1977_inst
    process(type_cast_1973_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1973_wire, type_cast_1976_wire_constant, tmp_var);
      ASHR_i32_i32_1977_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2060_inst
    process(type_cast_2056_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2056_wire, type_cast_2059_wire_constant, tmp_var);
      ASHR_i32_i32_2060_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2085_inst
    process(type_cast_2081_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2081_wire, type_cast_2084_wire_constant, tmp_var);
      ASHR_i32_i32_2085_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2393_inst
    process(type_cast_2389_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2389_wire, type_cast_2392_wire_constant, tmp_var);
      ASHR_i32_i32_2393_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2476_inst
    process(type_cast_2472_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2472_wire, type_cast_2475_wire_constant, tmp_var);
      ASHR_i32_i32_2476_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2501_inst
    process(type_cast_2497_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2497_wire, type_cast_2500_wire_constant, tmp_var);
      ASHR_i32_i32_2501_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2791_inst
    process(type_cast_2787_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2787_wire, type_cast_2790_wire_constant, tmp_var);
      ASHR_i32_i32_2791_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2874_inst
    process(type_cast_2870_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2870_wire, type_cast_2873_wire_constant, tmp_var);
      ASHR_i32_i32_2874_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2899_inst
    process(type_cast_2895_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2895_wire, type_cast_2898_wire_constant, tmp_var);
      ASHR_i32_i32_2899_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3195_inst
    process(type_cast_3191_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3191_wire, type_cast_3194_wire_constant, tmp_var);
      ASHR_i32_i32_3195_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3278_inst
    process(type_cast_3274_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3274_wire, type_cast_3277_wire_constant, tmp_var);
      ASHR_i32_i32_3278_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3303_inst
    process(type_cast_3299_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3299_wire, type_cast_3302_wire_constant, tmp_var);
      ASHR_i32_i32_3303_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3605_inst
    process(type_cast_3601_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3601_wire, type_cast_3604_wire_constant, tmp_var);
      ASHR_i32_i32_3605_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3688_inst
    process(type_cast_3684_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3684_wire, type_cast_3687_wire_constant, tmp_var);
      ASHR_i32_i32_3688_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3713_inst
    process(type_cast_3709_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3709_wire, type_cast_3712_wire_constant, tmp_var);
      ASHR_i32_i32_3713_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_555_inst
    process(type_cast_551_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_551_wire, type_cast_554_wire_constant, tmp_var);
      ASHR_i32_i32_555_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_617_inst
    process(type_cast_613_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_613_wire, type_cast_616_wire_constant, tmp_var);
      ASHR_i32_i32_617_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_755_inst
    process(type_cast_751_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_751_wire, type_cast_754_wire_constant, tmp_var);
      ASHR_i32_i32_755_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_839_inst
    process(type_cast_835_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_835_wire, type_cast_838_wire_constant, tmp_var);
      ASHR_i32_i32_839_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_864_inst
    process(type_cast_860_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_860_wire, type_cast_863_wire_constant, tmp_var);
      ASHR_i32_i32_864_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1341_inst
    process(conv436_1337, add442_1016) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv436_1337, add442_1016, tmp_var);
      cmp443_1342 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1366_inst
    process(conv451_1362, add458_1021) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv451_1362, add458_1021, tmp_var);
      cmp459_1367 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1755_inst
    process(conv653_1751, add660_1424) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv653_1751, add660_1424, tmp_var);
      cmp661_1756 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1781_inst
    process(conv669_1777, add676_1435) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv669_1777, add676_1435, tmp_var);
      cmp677_1782 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2153_inst
    process(conv874_2149, add880_1829) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv874_2149, add880_1829, tmp_var);
      cmp881_2154 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2178_inst
    process(conv889_2174, add896_1834) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv889_2174, add896_1834, tmp_var);
      cmp897_2179 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2569_inst
    process(conv1092_2565, add1099_2232) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1092_2565, add1099_2232, tmp_var);
      cmp1100_2570 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2595_inst
    process(conv1108_2591, add1116_2249) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1108_2591, add1116_2249, tmp_var);
      cmp1117_2596 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2967_inst
    process(conv1315_2963, add1321_2643) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1315_2963, add1321_2643, tmp_var);
      cmp1322_2968 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2992_inst
    process(conv1330_2988, add1338_2648) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1330_2988, add1338_2648, tmp_var);
      cmp1339_2993 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3371_inst
    process(conv1533_3367, add1540_3046) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1533_3367, add1540_3046, tmp_var);
      cmp1541_3372 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3397_inst
    process(conv1549_3393, add1555_3051) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1549_3393, add1555_3051, tmp_var);
      cmp1556_3398 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3781_inst
    process(conv1753_3777, add1759_3457) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1753_3777, add1759_3457, tmp_var);
      cmp1760_3782 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3806_inst
    process(conv1768_3802, add1774_3462) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv1768_3802, add1774_3462, tmp_var);
      cmp1775_3807 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_932_inst
    process(conv221_928, add228_574) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv221_928, add228_574, tmp_var);
      cmp229_933 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_958_inst
    process(conv237_954, add244_589) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv237_954, add244_589, tmp_var);
      cmp245_959 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_286_inst
    process(shr1839x_xmask_281) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr1839x_xmask_281, type_cast_285_wire_constant, tmp_var);
      cmp1840_287 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_499_inst
    process(indvarx_xnext_495, umax7_335) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_495, umax7_335, tmp_var);
      exitcond8_500 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1405_inst
    process(conv477_1400) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv477_1400, type_cast_1404_wire_constant, tmp_var);
      div478_1406 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2213_inst
    process(conv477_1400) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv477_1400, type_cast_2212_wire_constant, tmp_var);
      div916_2214 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3438_inst
    process(mul1579_3433) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1579_3433, type_cast_3437_wire_constant, tmp_var);
      div1580_3439 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_997_inst
    process(conv259_992) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv259_992, type_cast_996_wire_constant, tmp_var);
      div260_998 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1429_inst
    process(conv239_578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv239_578, type_cast_1428_wire_constant, tmp_var);
      div672_1430 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2243_inst
    process(mul1111_2238) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul1111_2238, type_cast_2242_wire_constant, tmp_var);
      div1112_2244 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_562_inst
    process(conv94_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv94_521, type_cast_561_wire_constant, tmp_var);
      div224_563 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_583_inst
    process(conv239_578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv239_578, type_cast_582_wire_constant, tmp_var);
      div240_584 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_321_inst
    process(tmp4_316) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_316, type_cast_320_wire_constant, tmp_var);
      tmp5_322 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3027_inst
    process(div478_1406) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(div478_1406, type_cast_3026_wire_constant, tmp_var);
      mul1359_3028 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3432_inst
    process(conv477_1400) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv477_1400, type_cast_3431_wire_constant, tmp_var);
      mul1579_3433 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1142_inst
    process(conv356_1138, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv356_1138, conv144_542, tmp_var);
      mul357_1143 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1147_inst
    process(conv315_1059, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv315_1059, conv150_557, tmp_var);
      mul363_1148 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1200_inst
    process(sub380_1196, conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub380_1196, conv92_517, tmp_var);
      mul381_1201 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1210_inst
    process(sub389_1206, conv171_619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub389_1206, conv171_619, tmp_var);
      mul390_1211 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1225_inst
    process(conv333_1096, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv333_1096, conv144_542, tmp_var);
      mul400_1226 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1230_inst
    process(conv315_1059, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv315_1059, conv150_557, tmp_var);
      mul406_1231 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1556_inst
    process(conv573_1552, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv573_1552, conv144_542, tmp_var);
      mul574_1557 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1561_inst
    process(conv531_1473, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv531_1473, conv150_557, tmp_var);
      mul580_1562 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1614_inst
    process(sub597_1610, conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub597_1610, conv92_517, tmp_var);
      mul598_1615 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1624_inst
    process(sub606_1620, conv171_619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub606_1620, conv171_619, tmp_var);
      mul607_1625 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1639_inst
    process(conv549_1510, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv549_1510, conv144_542, tmp_var);
      mul617_1640 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1644_inst
    process(conv531_1473, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv531_1473, conv150_557, tmp_var);
      mul623_1645 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1954_inst
    process(conv794_1950, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv794_1950, conv144_542, tmp_var);
      mul795_1955 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1959_inst
    process(conv753_1871, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv753_1871, conv150_557, tmp_var);
      mul801_1960 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2012_inst
    process(sub818_2008, conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub818_2008, conv92_517, tmp_var);
      mul819_2013 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2022_inst
    process(sub827_2018, conv171_619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub827_2018, conv171_619, tmp_var);
      mul828_2023 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2037_inst
    process(conv771_1908, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv771_1908, conv144_542, tmp_var);
      mul838_2038 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2042_inst
    process(conv753_1871, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv753_1871, conv150_557, tmp_var);
      mul844_2043 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2237_inst
    process(conv239_578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv239_578, type_cast_2236_wire_constant, tmp_var);
      mul1111_2238 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2370_inst
    process(conv1012_2366, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1012_2366, conv144_542, tmp_var);
      mul1013_2371 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2375_inst
    process(conv969_2287, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv969_2287, conv150_557, tmp_var);
      mul1019_2376 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2428_inst
    process(sub1036_2424, conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1036_2424, conv92_517, tmp_var);
      mul1037_2429 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2438_inst
    process(sub1045_2434, conv171_619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1045_2434, conv171_619, tmp_var);
      mul1046_2439 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2453_inst
    process(conv988_2324, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv988_2324, conv144_542, tmp_var);
      mul1056_2454 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2458_inst
    process(conv969_2287, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv969_2287, conv150_557, tmp_var);
      mul1062_2459 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2768_inst
    process(conv1235_2764, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1235_2764, conv144_542, tmp_var);
      mul1236_2769 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2773_inst
    process(conv1193_2685, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1193_2685, conv150_557, tmp_var);
      mul1242_2774 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2826_inst
    process(sub1259_2822, conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1259_2822, conv92_517, tmp_var);
      mul1260_2827 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2836_inst
    process(sub1268_2832, conv171_619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1268_2832, conv171_619, tmp_var);
      mul1269_2837 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2851_inst
    process(conv1212_2722, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1212_2722, conv144_542, tmp_var);
      mul1279_2852 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2856_inst
    process(conv1193_2685, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1193_2685, conv150_557, tmp_var);
      mul1285_2857 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3172_inst
    process(conv1453_3168, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1453_3168, conv144_542, tmp_var);
      mul1454_3173 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3177_inst
    process(conv1412_3089, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1412_3089, conv150_557, tmp_var);
      mul1460_3178 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3230_inst
    process(sub1477_3226, conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1477_3226, conv92_517, tmp_var);
      mul1478_3231 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3240_inst
    process(sub1486_3236, conv171_619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1486_3236, conv171_619, tmp_var);
      mul1487_3241 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3255_inst
    process(conv1429_3126, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1429_3126, conv144_542, tmp_var);
      mul1497_3256 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3260_inst
    process(conv1412_3089, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1412_3089, conv150_557, tmp_var);
      mul1503_3261 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3582_inst
    process(conv1673_3578, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1673_3578, conv144_542, tmp_var);
      mul1674_3583 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3587_inst
    process(conv1633_3499, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1633_3499, conv150_557, tmp_var);
      mul1680_3588 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3640_inst
    process(sub1697_3636, conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1697_3636, conv92_517, tmp_var);
      mul1698_3641 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3650_inst
    process(sub1706_3646, conv171_619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub1706_3646, conv171_619, tmp_var);
      mul1707_3651 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3665_inst
    process(conv1650_3536, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1650_3536, conv144_542, tmp_var);
      mul1717_3666 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3670_inst
    process(conv1633_3499, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1633_3499, conv150_557, tmp_var);
      mul1723_3671 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3849_inst
    process(conv1790_3845, conv1788_3841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv1790_3845, conv1788_3841, tmp_var);
      mul1791_3850 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3854_inst
    process(mul1791_3850, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul1791_3850, conv144_542, tmp_var);
      mul1794_3855 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_533_inst
    process(conv99_525, conv101_529) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv99_525, conv101_529, tmp_var);
      mul102_534 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_609_inst
    process(mul95_605, conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul95_605, conv92_517, tmp_var);
      sext_610 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_732_inst
    process(conv146_728, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv146_728, conv144_542, tmp_var);
      mul147_733 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_737_inst
    process(conv108_649, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv108_649, conv150_557, tmp_var);
      mul153_738 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_791_inst
    process(sub_787, conv92_517) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub_787, conv92_517, tmp_var);
      mul168_792 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_801_inst
    process(sub176_797, conv171_619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub176_797, conv171_619, tmp_var);
      mul177_802 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_816_inst
    process(conv124_686, conv144_542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv124_686, conv144_542, tmp_var);
      mul187_817 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_821_inst
    process(conv108_649, conv150_557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv108_649, conv150_557, tmp_var);
      mul193_822 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_269_inst
    process(conv10_261, conv_257) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv10_261, conv_257, tmp_var);
      mul_270 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_274_inst
    process(mul_270, conv12_265) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_270, conv12_265, tmp_var);
      mul13_275 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_306_inst
    process(tmp_298, tmp1_302) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_298, tmp1_302, tmp_var);
      tmp2_307 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_315_inst
    process(tmp2_307, tmp3_311) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_307, tmp3_311, tmp_var);
      tmp4_316 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_376_inst
    process(shl_365, conv25_372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_365, conv25_372, tmp_var);
      add_377 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_394_inst
    process(shl27_383, conv30_390) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_383, conv30_390, tmp_var);
      add31_395 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_412_inst
    process(shl33_401, conv36_408) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl33_401, conv36_408, tmp_var);
      add37_413 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_430_inst
    process(shl39_419, conv42_426) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl39_419, conv42_426, tmp_var);
      add43_431 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_448_inst
    process(shl45_437, conv48_444) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_437, conv48_444, tmp_var);
      add49_449 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_466_inst
    process(shl51_455, conv54_462) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl51_455, conv54_462, tmp_var);
      add55_467 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_484_inst
    process(shl57_473, conv60_480) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl57_473, conv60_480, tmp_var);
      add61_485 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1010_inst
    process(conv317_1005) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv317_1005, type_cast_1009_wire_constant, tmp_var);
      shl441_1011 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1418_inst
    process(conv533_1413) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv533_1413, type_cast_1417_wire_constant, tmp_var);
      shl659_1419 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1823_inst
    process(conv755_1818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv755_1818, type_cast_1822_wire_constant, tmp_var);
      shl879_1824 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2226_inst
    process(conv971_2221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv971_2221, type_cast_2225_wire_constant, tmp_var);
      shl1098_2227 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2637_inst
    process(conv1195_2632) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1195_2632, type_cast_2636_wire_constant, tmp_var);
      shl1320_2638 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3040_inst
    process(conv1414_3035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1414_3035, type_cast_3039_wire_constant, tmp_var);
      shl1539_3041 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3451_inst
    process(conv1635_3446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1635_3446, type_cast_3450_wire_constant, tmp_var);
      shl1758_3452 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_547_inst
    process(mul102_534) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul102_534, type_cast_546_wire_constant, tmp_var);
      sext1848_548 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_568_inst
    process(conv110_538) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv110_538, type_cast_567_wire_constant, tmp_var);
      shl227_569 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_604_inst
    process(conv94_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv94_521, type_cast_603_wire_constant, tmp_var);
      mul95_605 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_364_inst
    process(conv21_359) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv21_359, type_cast_363_wire_constant, tmp_var);
      shl_365 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_382_inst
    process(add_377) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_377, type_cast_381_wire_constant, tmp_var);
      shl27_383 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_400_inst
    process(add31_395) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add31_395, type_cast_399_wire_constant, tmp_var);
      shl33_401 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_418_inst
    process(add37_413) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add37_413, type_cast_417_wire_constant, tmp_var);
      shl39_419 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_436_inst
    process(add43_431) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add43_431, type_cast_435_wire_constant, tmp_var);
      shl45_437 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_454_inst
    process(add49_449) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add49_449, type_cast_453_wire_constant, tmp_var);
      shl51_455 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_472_inst
    process(add55_467) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add55_467, type_cast_471_wire_constant, tmp_var);
      shl57_473 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1065_inst
    process(type_cast_1062_wire, type_cast_1064_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1062_wire, type_cast_1064_wire, tmp_var);
      cmp318_1066 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1078_inst
    process(type_cast_1075_wire, type_cast_1077_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1075_wire, type_cast_1077_wire, tmp_var);
      cmp329_1079 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1102_inst
    process(type_cast_1099_wire, type_cast_1101_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1099_wire, type_cast_1101_wire, tmp_var);
      cmp336_1103 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1115_inst
    process(type_cast_1112_wire, type_cast_1114_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1112_wire, type_cast_1114_wire, tmp_var);
      cmp346_1116 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1310_inst
    process(type_cast_1307_wire, type_cast_1309_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1307_wire, type_cast_1309_wire, tmp_var);
      cmp425_1311 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1479_inst
    process(type_cast_1476_wire, type_cast_1478_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1476_wire, type_cast_1478_wire, tmp_var);
      cmp534_1480 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1492_inst
    process(type_cast_1489_wire, type_cast_1491_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1489_wire, type_cast_1491_wire, tmp_var);
      cmp545_1493 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1516_inst
    process(type_cast_1513_wire, type_cast_1515_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1513_wire, type_cast_1515_wire, tmp_var);
      cmp552_1517 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1529_inst
    process(type_cast_1526_wire, type_cast_1528_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1526_wire, type_cast_1528_wire, tmp_var);
      cmp563_1530 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1724_inst
    process(type_cast_1721_wire, type_cast_1723_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1721_wire, type_cast_1723_wire, tmp_var);
      cmp642_1725 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1877_inst
    process(type_cast_1874_wire, type_cast_1876_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1874_wire, type_cast_1876_wire, tmp_var);
      cmp756_1878 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1890_inst
    process(type_cast_1887_wire, type_cast_1889_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1887_wire, type_cast_1889_wire, tmp_var);
      cmp767_1891 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1914_inst
    process(type_cast_1911_wire, type_cast_1913_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1911_wire, type_cast_1913_wire, tmp_var);
      cmp774_1915 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1927_inst
    process(type_cast_1924_wire, type_cast_1926_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1924_wire, type_cast_1926_wire, tmp_var);
      cmp784_1928 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2122_inst
    process(type_cast_2119_wire, type_cast_2121_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2119_wire, type_cast_2121_wire, tmp_var);
      cmp863_2123 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2293_inst
    process(type_cast_2290_wire, type_cast_2292_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2290_wire, type_cast_2292_wire, tmp_var);
      cmp972_2294 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2306_inst
    process(type_cast_2303_wire, type_cast_2305_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2303_wire, type_cast_2305_wire, tmp_var);
      cmp984_2307 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2330_inst
    process(type_cast_2327_wire, type_cast_2329_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2327_wire, type_cast_2329_wire, tmp_var);
      cmp991_2331 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2343_inst
    process(type_cast_2340_wire, type_cast_2342_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2340_wire, type_cast_2342_wire, tmp_var);
      cmp1002_2344 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2538_inst
    process(type_cast_2535_wire, type_cast_2537_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2535_wire, type_cast_2537_wire, tmp_var);
      cmp1081_2539 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2691_inst
    process(type_cast_2688_wire, type_cast_2690_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2688_wire, type_cast_2690_wire, tmp_var);
      cmp1196_2692 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2704_inst
    process(type_cast_2701_wire, type_cast_2703_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2701_wire, type_cast_2703_wire, tmp_var);
      cmp1208_2705 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2728_inst
    process(type_cast_2725_wire, type_cast_2727_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2725_wire, type_cast_2727_wire, tmp_var);
      cmp1215_2729 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2741_inst
    process(type_cast_2738_wire, type_cast_2740_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2738_wire, type_cast_2740_wire, tmp_var);
      cmp1225_2742 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_2936_inst
    process(type_cast_2933_wire, type_cast_2935_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_2933_wire, type_cast_2935_wire, tmp_var);
      cmp1304_2937 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3095_inst
    process(type_cast_3092_wire, type_cast_3094_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3092_wire, type_cast_3094_wire, tmp_var);
      cmp1415_3096 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3108_inst
    process(type_cast_3105_wire, type_cast_3107_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3105_wire, type_cast_3107_wire, tmp_var);
      cmp1425_3109 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3132_inst
    process(type_cast_3129_wire, type_cast_3131_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3129_wire, type_cast_3131_wire, tmp_var);
      cmp1432_3133 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3145_inst
    process(type_cast_3142_wire, type_cast_3144_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3142_wire, type_cast_3144_wire, tmp_var);
      cmp1443_3146 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3340_inst
    process(type_cast_3337_wire, type_cast_3339_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3337_wire, type_cast_3339_wire, tmp_var);
      cmp1522_3341 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3505_inst
    process(type_cast_3502_wire, type_cast_3504_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3502_wire, type_cast_3504_wire, tmp_var);
      cmp1636_3506 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3518_inst
    process(type_cast_3515_wire, type_cast_3517_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3515_wire, type_cast_3517_wire, tmp_var);
      cmp1646_3519 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3542_inst
    process(type_cast_3539_wire, type_cast_3541_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3539_wire, type_cast_3541_wire, tmp_var);
      cmp1653_3543 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3555_inst
    process(type_cast_3552_wire, type_cast_3554_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3552_wire, type_cast_3554_wire, tmp_var);
      cmp1663_3556 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_3750_inst
    process(type_cast_3747_wire, type_cast_3749_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_3747_wire, type_cast_3749_wire, tmp_var);
      cmp1742_3751 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_655_inst
    process(type_cast_652_wire, type_cast_654_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_652_wire, type_cast_654_wire, tmp_var);
      cmp111_656 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_668_inst
    process(type_cast_665_wire, type_cast_667_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_665_wire, type_cast_667_wire, tmp_var);
      cmp120_669 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_692_inst
    process(type_cast_689_wire, type_cast_691_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_689_wire, type_cast_691_wire, tmp_var);
      cmp127_693 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_705_inst
    process(type_cast_702_wire, type_cast_704_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_702_wire, type_cast_704_wire, tmp_var);
      cmp138_706 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_901_inst
    process(type_cast_898_wire, type_cast_900_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_898_wire, type_cast_900_wire, tmp_var);
      cmp210_902 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1195_inst
    process(conv333_1096, conv317_1005) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv333_1096, conv317_1005, tmp_var);
      sub380_1196 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1205_inst
    process(conv315_1059, conv317_1005) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv315_1059, conv317_1005, tmp_var);
      sub389_1206 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1609_inst
    process(conv549_1510, conv533_1413) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv549_1510, conv533_1413, tmp_var);
      sub597_1610 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1619_inst
    process(conv531_1473, conv533_1413) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv531_1473, conv533_1413, tmp_var);
      sub606_1620 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2007_inst
    process(conv771_1908, conv755_1818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv771_1908, conv755_1818, tmp_var);
      sub818_2008 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2017_inst
    process(conv753_1871, conv755_1818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv753_1871, conv755_1818, tmp_var);
      sub827_2018 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2423_inst
    process(conv988_2324, conv971_2221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv988_2324, conv971_2221, tmp_var);
      sub1036_2424 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2433_inst
    process(conv969_2287, conv971_2221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv969_2287, conv971_2221, tmp_var);
      sub1045_2434 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2821_inst
    process(conv1212_2722, conv1195_2632) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1212_2722, conv1195_2632, tmp_var);
      sub1259_2822 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2831_inst
    process(conv1193_2685, conv1195_2632) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1193_2685, conv1195_2632, tmp_var);
      sub1268_2832 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3225_inst
    process(conv1429_3126, conv1414_3035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1429_3126, conv1414_3035, tmp_var);
      sub1477_3226 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3235_inst
    process(conv1412_3089, conv1414_3035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1412_3089, conv1414_3035, tmp_var);
      sub1486_3236 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3635_inst
    process(conv1650_3536, conv1635_3446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1650_3536, conv1635_3446, tmp_var);
      sub1697_3636 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_3645_inst
    process(conv1633_3499, conv1635_3446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv1633_3499, conv1635_3446, tmp_var);
      sub1706_3646 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_786_inst
    process(conv124_686, conv110_538) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv124_686, conv110_538, tmp_var);
      sub_787 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_796_inst
    process(conv108_649, conv110_538) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv108_649, conv110_538, tmp_var);
      sub176_797 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_327_inst
    process(tmp5_322) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp5_322, type_cast_326_wire_constant, tmp_var);
      tmp6_328 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1071_inst
    process(cmp318_1066) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp318_1066, type_cast_1070_wire_constant, tmp_var);
      cmp318x_xnot_1072 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1108_inst
    process(cmp336_1103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp336_1103, type_cast_1107_wire_constant, tmp_var);
      cmp336x_xnot_1109 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1485_inst
    process(cmp534_1480) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp534_1480, type_cast_1484_wire_constant, tmp_var);
      cmp534x_xnot_1486 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1522_inst
    process(cmp552_1517) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp552_1517, type_cast_1521_wire_constant, tmp_var);
      cmp552x_xnot_1523 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1883_inst
    process(cmp756_1878) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp756_1878, type_cast_1882_wire_constant, tmp_var);
      cmp756x_xnot_1884 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1920_inst
    process(cmp774_1915) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp774_1915, type_cast_1919_wire_constant, tmp_var);
      cmp774x_xnot_1921 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_2299_inst
    process(cmp972_2294) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp972_2294, type_cast_2298_wire_constant, tmp_var);
      cmp972x_xnot_2300 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_2336_inst
    process(cmp991_2331) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp991_2331, type_cast_2335_wire_constant, tmp_var);
      cmp991x_xnot_2337 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_2697_inst
    process(cmp1196_2692) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp1196_2692, type_cast_2696_wire_constant, tmp_var);
      cmp1196x_xnot_2698 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_2734_inst
    process(cmp1215_2729) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp1215_2729, type_cast_2733_wire_constant, tmp_var);
      cmp1215x_xnot_2735 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_3101_inst
    process(cmp1415_3096) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp1415_3096, type_cast_3100_wire_constant, tmp_var);
      cmp1415x_xnot_3102 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_3138_inst
    process(cmp1432_3133) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp1432_3133, type_cast_3137_wire_constant, tmp_var);
      cmp1432x_xnot_3139 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_3511_inst
    process(cmp1636_3506) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp1636_3506, type_cast_3510_wire_constant, tmp_var);
      cmp1636x_xnot_3512 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_3548_inst
    process(cmp1653_3543) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp1653_3543, type_cast_3547_wire_constant, tmp_var);
      cmp1653x_xnot_3549 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_661_inst
    process(cmp111_656) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp111_656, type_cast_660_wire_constant, tmp_var);
      cmp111x_xnot_662 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_698_inst
    process(cmp127_693) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp127_693, type_cast_697_wire_constant, tmp_var);
      cmp127x_xnot_699 <= tmp_var; --
    end process;
    -- shared split operator group (339) : array_obj_ref_1177_index_offset 
    ApIntAdd_group_339: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom367_1176_scaled;
      array_obj_ref_1177_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1177_index_offset_req_0;
      array_obj_ref_1177_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1177_index_offset_req_1;
      array_obj_ref_1177_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_339_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_339_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_339",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 339
    -- shared split operator group (340) : array_obj_ref_1260_index_offset 
    ApIntAdd_group_340: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom410_1259_scaled;
      array_obj_ref_1260_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1260_index_offset_req_0;
      array_obj_ref_1260_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1260_index_offset_req_1;
      array_obj_ref_1260_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_340_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_340_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_340",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 340
    -- shared split operator group (341) : array_obj_ref_1285_index_offset 
    ApIntAdd_group_341: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom415_1284_scaled;
      array_obj_ref_1285_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1285_index_offset_req_0;
      array_obj_ref_1285_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1285_index_offset_req_1;
      array_obj_ref_1285_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_341_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_341_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_341",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 341
    -- shared split operator group (342) : array_obj_ref_1591_index_offset 
    ApIntAdd_group_342: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom584_1590_scaled;
      array_obj_ref_1591_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1591_index_offset_req_0;
      array_obj_ref_1591_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1591_index_offset_req_1;
      array_obj_ref_1591_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_342_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_342_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_342",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 342
    -- shared split operator group (343) : array_obj_ref_1674_index_offset 
    ApIntAdd_group_343: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom627_1673_scaled;
      array_obj_ref_1674_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1674_index_offset_req_0;
      array_obj_ref_1674_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1674_index_offset_req_1;
      array_obj_ref_1674_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_343_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_343_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_343",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 343
    -- shared split operator group (344) : array_obj_ref_1699_index_offset 
    ApIntAdd_group_344: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom632_1698_scaled;
      array_obj_ref_1699_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1699_index_offset_req_0;
      array_obj_ref_1699_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1699_index_offset_req_1;
      array_obj_ref_1699_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_344_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_344_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_344",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 344
    -- shared split operator group (345) : array_obj_ref_1989_index_offset 
    ApIntAdd_group_345: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom805_1988_scaled;
      array_obj_ref_1989_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1989_index_offset_req_0;
      array_obj_ref_1989_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1989_index_offset_req_1;
      array_obj_ref_1989_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_345_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_345_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_345",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 345
    -- shared split operator group (346) : array_obj_ref_2072_index_offset 
    ApIntAdd_group_346: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom848_2071_scaled;
      array_obj_ref_2072_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2072_index_offset_req_0;
      array_obj_ref_2072_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2072_index_offset_req_1;
      array_obj_ref_2072_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_346_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_346_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_346",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 346
    -- shared split operator group (347) : array_obj_ref_2097_index_offset 
    ApIntAdd_group_347: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom853_2096_scaled;
      array_obj_ref_2097_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2097_index_offset_req_0;
      array_obj_ref_2097_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2097_index_offset_req_1;
      array_obj_ref_2097_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_347_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_347_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_347",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 347
    -- shared split operator group (348) : array_obj_ref_2405_index_offset 
    ApIntAdd_group_348: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1023_2404_scaled;
      array_obj_ref_2405_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2405_index_offset_req_0;
      array_obj_ref_2405_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2405_index_offset_req_1;
      array_obj_ref_2405_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_348_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_348_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_348",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 348
    -- shared split operator group (349) : array_obj_ref_2488_index_offset 
    ApIntAdd_group_349: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1066_2487_scaled;
      array_obj_ref_2488_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2488_index_offset_req_0;
      array_obj_ref_2488_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2488_index_offset_req_1;
      array_obj_ref_2488_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_349_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_349_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_349",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 349
    -- shared split operator group (350) : array_obj_ref_2513_index_offset 
    ApIntAdd_group_350: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1071_2512_scaled;
      array_obj_ref_2513_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2513_index_offset_req_0;
      array_obj_ref_2513_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2513_index_offset_req_1;
      array_obj_ref_2513_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_350_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_350_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_350",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 350
    -- shared split operator group (351) : array_obj_ref_2803_index_offset 
    ApIntAdd_group_351: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1246_2802_scaled;
      array_obj_ref_2803_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2803_index_offset_req_0;
      array_obj_ref_2803_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2803_index_offset_req_1;
      array_obj_ref_2803_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_351_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_351_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_351",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 351
    -- shared split operator group (352) : array_obj_ref_2886_index_offset 
    ApIntAdd_group_352: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1289_2885_scaled;
      array_obj_ref_2886_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2886_index_offset_req_0;
      array_obj_ref_2886_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2886_index_offset_req_1;
      array_obj_ref_2886_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_352_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_352_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_352",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 352
    -- shared split operator group (353) : array_obj_ref_2911_index_offset 
    ApIntAdd_group_353: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1294_2910_scaled;
      array_obj_ref_2911_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2911_index_offset_req_0;
      array_obj_ref_2911_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2911_index_offset_req_1;
      array_obj_ref_2911_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_353_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_353_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_353",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 353
    -- shared split operator group (354) : array_obj_ref_3207_index_offset 
    ApIntAdd_group_354: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1464_3206_scaled;
      array_obj_ref_3207_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3207_index_offset_req_0;
      array_obj_ref_3207_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3207_index_offset_req_1;
      array_obj_ref_3207_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_354_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_354_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_354",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 354
    -- shared split operator group (355) : array_obj_ref_3290_index_offset 
    ApIntAdd_group_355: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1507_3289_scaled;
      array_obj_ref_3290_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3290_index_offset_req_0;
      array_obj_ref_3290_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3290_index_offset_req_1;
      array_obj_ref_3290_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_355_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_355_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_355",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 355
    -- shared split operator group (356) : array_obj_ref_3315_index_offset 
    ApIntAdd_group_356: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1512_3314_scaled;
      array_obj_ref_3315_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3315_index_offset_req_0;
      array_obj_ref_3315_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3315_index_offset_req_1;
      array_obj_ref_3315_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_356_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_356_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_356",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 356
    -- shared split operator group (357) : array_obj_ref_350_index_offset 
    ApIntAdd_group_357: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_349_scaled;
      array_obj_ref_350_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_350_index_offset_req_0;
      array_obj_ref_350_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_350_index_offset_req_1;
      array_obj_ref_350_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_357_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_357_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_357",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 357
    -- shared split operator group (358) : array_obj_ref_3617_index_offset 
    ApIntAdd_group_358: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1684_3616_scaled;
      array_obj_ref_3617_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3617_index_offset_req_0;
      array_obj_ref_3617_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3617_index_offset_req_1;
      array_obj_ref_3617_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_358_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_358_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_358",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 358
    -- shared split operator group (359) : array_obj_ref_3700_index_offset 
    ApIntAdd_group_359: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1727_3699_scaled;
      array_obj_ref_3700_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3700_index_offset_req_0;
      array_obj_ref_3700_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3700_index_offset_req_1;
      array_obj_ref_3700_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_359_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_359_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_359",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 359
    -- shared split operator group (360) : array_obj_ref_3725_index_offset 
    ApIntAdd_group_360: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom1732_3724_scaled;
      array_obj_ref_3725_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3725_index_offset_req_0;
      array_obj_ref_3725_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3725_index_offset_req_1;
      array_obj_ref_3725_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_360_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_360_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_360",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 360
    -- shared split operator group (361) : array_obj_ref_768_index_offset 
    ApIntAdd_group_361: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom157_767_scaled;
      array_obj_ref_768_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_768_index_offset_req_0;
      array_obj_ref_768_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_768_index_offset_req_1;
      array_obj_ref_768_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_361_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_361_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_361",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 361
    -- shared split operator group (362) : array_obj_ref_851_index_offset 
    ApIntAdd_group_362: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom197_850_scaled;
      array_obj_ref_851_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_851_index_offset_req_0;
      array_obj_ref_851_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_851_index_offset_req_1;
      array_obj_ref_851_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_362_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_362_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_362",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 362
    -- shared split operator group (363) : array_obj_ref_876_index_offset 
    ApIntAdd_group_363: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom202_875_scaled;
      array_obj_ref_876_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_876_index_offset_req_0;
      array_obj_ref_876_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_876_index_offset_req_1;
      array_obj_ref_876_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_363_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_363_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_363",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 363
    -- unary operator type_cast_1057_inst
    process(i263x_x2_1040) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i263x_x2_1040, tmp_var);
      type_cast_1057_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1094_inst
    process(j309x_x1_1034) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j309x_x1_1034, tmp_var);
      type_cast_1094_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1131_inst
    process(k255x_x1_1047) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k255x_x1_1047, tmp_var);
      type_cast_1131_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1136_inst
    process(j309x_x1_1034) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j309x_x1_1034, tmp_var);
      type_cast_1136_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1170_inst
    process(shr366_1167) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr366_1167, tmp_var);
      type_cast_1170_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1189_inst
    process(k255x_x1_1047) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k255x_x1_1047, tmp_var);
      type_cast_1189_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1253_inst
    process(shr409_1250) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr409_1250, tmp_var);
      type_cast_1253_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1278_inst
    process(shr414_1275) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr414_1275, tmp_var);
      type_cast_1278_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1296_inst
    process(k255x_x1_1047) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k255x_x1_1047, tmp_var);
      type_cast_1296_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1335_inst
    process(inc434_1332) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc434_1332, tmp_var);
      type_cast_1335_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1360_inst
    process(inc448x_xi263x_x2_1351) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc448x_xi263x_x2_1351, tmp_var);
      type_cast_1360_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1471_inst
    process(i475x_x2_1455) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i475x_x2_1455, tmp_var);
      type_cast_1471_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1508_inst
    process(j525x_x1_1461) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j525x_x1_1461, tmp_var);
      type_cast_1508_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1545_inst
    process(k471x_x1_1448) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k471x_x1_1448, tmp_var);
      type_cast_1545_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1550_inst
    process(j525x_x1_1461) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j525x_x1_1461, tmp_var);
      type_cast_1550_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1584_inst
    process(shr583_1581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr583_1581, tmp_var);
      type_cast_1584_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1603_inst
    process(k471x_x1_1448) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k471x_x1_1448, tmp_var);
      type_cast_1603_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1667_inst
    process(shr626_1664) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr626_1664, tmp_var);
      type_cast_1667_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1692_inst
    process(shr631_1689) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr631_1689, tmp_var);
      type_cast_1692_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1710_inst
    process(k471x_x1_1448) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k471x_x1_1448, tmp_var);
      type_cast_1710_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1749_inst
    process(inc651_1746) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc651_1746, tmp_var);
      type_cast_1749_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1775_inst
    process(inc666x_xi475x_x2_1765) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc666x_xi475x_x2_1765, tmp_var);
      type_cast_1775_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1869_inst
    process(i697x_x2_1854) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i697x_x2_1854, tmp_var);
      type_cast_1869_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1906_inst
    process(j747x_x1_1860) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j747x_x1_1860, tmp_var);
      type_cast_1906_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1943_inst
    process(k689x_x1_1847) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k689x_x1_1847, tmp_var);
      type_cast_1943_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1948_inst
    process(j747x_x1_1860) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j747x_x1_1860, tmp_var);
      type_cast_1948_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1982_inst
    process(shr804_1979) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr804_1979, tmp_var);
      type_cast_1982_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2001_inst
    process(k689x_x1_1847) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k689x_x1_1847, tmp_var);
      type_cast_2001_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2065_inst
    process(shr847_2062) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr847_2062, tmp_var);
      type_cast_2065_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2090_inst
    process(shr852_2087) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr852_2087, tmp_var);
      type_cast_2090_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2108_inst
    process(k689x_x1_1847) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k689x_x1_1847, tmp_var);
      type_cast_2108_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2147_inst
    process(inc872_2144) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc872_2144, tmp_var);
      type_cast_2147_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2172_inst
    process(inc886x_xi697x_x2_2163) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc886x_xi697x_x2_2163, tmp_var);
      type_cast_2172_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2285_inst
    process(i913x_x2_2269) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i913x_x2_2269, tmp_var);
      type_cast_2285_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2322_inst
    process(j963x_x1_2275) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j963x_x1_2275, tmp_var);
      type_cast_2322_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2359_inst
    process(k909x_x1_2262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k909x_x1_2262, tmp_var);
      type_cast_2359_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2364_inst
    process(j963x_x1_2275) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j963x_x1_2275, tmp_var);
      type_cast_2364_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2398_inst
    process(shr1022_2395) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1022_2395, tmp_var);
      type_cast_2398_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2417_inst
    process(k909x_x1_2262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k909x_x1_2262, tmp_var);
      type_cast_2417_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2481_inst
    process(shr1065_2478) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1065_2478, tmp_var);
      type_cast_2481_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2506_inst
    process(shr1070_2503) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1070_2503, tmp_var);
      type_cast_2506_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2524_inst
    process(k909x_x1_2262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k909x_x1_2262, tmp_var);
      type_cast_2524_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2563_inst
    process(inc1090_2560) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1090_2560, tmp_var);
      type_cast_2563_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2589_inst
    process(inc1105x_xi913x_x2_2579) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1105x_xi913x_x2_2579, tmp_var);
      type_cast_2589_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2683_inst
    process(i1137x_x2_2668) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1137x_x2_2668, tmp_var);
      type_cast_2683_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2720_inst
    process(j1187x_x1_2674) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1187x_x1_2674, tmp_var);
      type_cast_2720_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2757_inst
    process(k1129x_x1_2661) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1129x_x1_2661, tmp_var);
      type_cast_2757_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2762_inst
    process(j1187x_x1_2674) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1187x_x1_2674, tmp_var);
      type_cast_2762_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2796_inst
    process(shr1245_2793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1245_2793, tmp_var);
      type_cast_2796_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2815_inst
    process(k1129x_x1_2661) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1129x_x1_2661, tmp_var);
      type_cast_2815_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2879_inst
    process(shr1288_2876) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1288_2876, tmp_var);
      type_cast_2879_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2904_inst
    process(shr1293_2901) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1293_2901, tmp_var);
      type_cast_2904_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2922_inst
    process(k1129x_x1_2661) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1129x_x1_2661, tmp_var);
      type_cast_2922_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2961_inst
    process(inc1313_2958) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1313_2958, tmp_var);
      type_cast_2961_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2986_inst
    process(inc1327x_xi1137x_x2_2977) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1327x_xi1137x_x2_2977, tmp_var);
      type_cast_2986_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3087_inst
    process(i1355x_x2_3071) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1355x_x2_3071, tmp_var);
      type_cast_3087_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3124_inst
    process(j1406x_x1_3077) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1406x_x1_3077, tmp_var);
      type_cast_3124_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3161_inst
    process(k1351x_x1_3064) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1351x_x1_3064, tmp_var);
      type_cast_3161_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3166_inst
    process(j1406x_x1_3077) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1406x_x1_3077, tmp_var);
      type_cast_3166_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3200_inst
    process(shr1463_3197) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1463_3197, tmp_var);
      type_cast_3200_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3219_inst
    process(k1351x_x1_3064) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1351x_x1_3064, tmp_var);
      type_cast_3219_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3283_inst
    process(shr1506_3280) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1506_3280, tmp_var);
      type_cast_3283_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3308_inst
    process(shr1511_3305) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1511_3305, tmp_var);
      type_cast_3308_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3326_inst
    process(k1351x_x1_3064) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1351x_x1_3064, tmp_var);
      type_cast_3326_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3365_inst
    process(inc1531_3362) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1531_3362, tmp_var);
      type_cast_3365_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3391_inst
    process(inc1546x_xi1355x_x2_3381) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1546x_xi1355x_x2_3381, tmp_var);
      type_cast_3391_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3497_inst
    process(i1576x_x2_3482) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i1576x_x2_3482, tmp_var);
      type_cast_3497_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3534_inst
    process(j1627x_x1_3488) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1627x_x1_3488, tmp_var);
      type_cast_3534_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3571_inst
    process(k1568x_x1_3475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1568x_x1_3475, tmp_var);
      type_cast_3571_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3576_inst
    process(j1627x_x1_3488) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", j1627x_x1_3488, tmp_var);
      type_cast_3576_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3610_inst
    process(shr1683_3607) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1683_3607, tmp_var);
      type_cast_3610_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3629_inst
    process(k1568x_x1_3475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1568x_x1_3475, tmp_var);
      type_cast_3629_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3693_inst
    process(shr1726_3690) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1726_3690, tmp_var);
      type_cast_3693_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3718_inst
    process(shr1731_3715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr1731_3715, tmp_var);
      type_cast_3718_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3736_inst
    process(k1568x_x1_3475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", k1568x_x1_3475, tmp_var);
      type_cast_3736_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3775_inst
    process(inc1751_3772) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1751_3772, tmp_var);
      type_cast_3775_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3800_inst
    process(inc1765x_xi1576x_x2_3791) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc1765x_xi1576x_x2_3791, tmp_var);
      type_cast_3800_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_647_inst
    process(i68x_x2_630) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", i68x_x2_630, tmp_var);
      type_cast_647_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_684_inst
    process(jx_x1_622) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_622, tmp_var);
      type_cast_684_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_721_inst
    process(kx_x1_637) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_637, tmp_var);
      type_cast_721_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_726_inst
    process(jx_x1_622) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", jx_x1_622, tmp_var);
      type_cast_726_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_761_inst
    process(shr156_757) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr156_757, tmp_var);
      type_cast_761_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_780_inst
    process(kx_x1_637) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_637, tmp_var);
      type_cast_780_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_844_inst
    process(shr196_841) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr196_841, tmp_var);
      type_cast_844_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_869_inst
    process(shr201_866) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr201_866, tmp_var);
      type_cast_869_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_887_inst
    process(kx_x1_637) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", kx_x1_637, tmp_var);
      type_cast_887_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_926_inst
    process(inc219_923) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc219_923, tmp_var);
      type_cast_926_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_952_inst
    process(inc234x_xi68x_x2_942) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc234x_xi68x_x2_942, tmp_var);
      type_cast_952_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_pad_1000_load_0 LOAD_pad_512_load_0 LOAD_pad_3441_load_0 LOAD_pad_1408_load_0 LOAD_pad_1813_load_0 LOAD_pad_2216_load_0 LOAD_pad_2627_load_0 LOAD_pad_3030_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= LOAD_pad_1000_load_0_req_0;
      reqL_unguarded(6) <= LOAD_pad_512_load_0_req_0;
      reqL_unguarded(5) <= LOAD_pad_3441_load_0_req_0;
      reqL_unguarded(4) <= LOAD_pad_1408_load_0_req_0;
      reqL_unguarded(3) <= LOAD_pad_1813_load_0_req_0;
      reqL_unguarded(2) <= LOAD_pad_2216_load_0_req_0;
      reqL_unguarded(1) <= LOAD_pad_2627_load_0_req_0;
      reqL_unguarded(0) <= LOAD_pad_3030_load_0_req_0;
      LOAD_pad_1000_load_0_ack_0 <= ackL_unguarded(7);
      LOAD_pad_512_load_0_ack_0 <= ackL_unguarded(6);
      LOAD_pad_3441_load_0_ack_0 <= ackL_unguarded(5);
      LOAD_pad_1408_load_0_ack_0 <= ackL_unguarded(4);
      LOAD_pad_1813_load_0_ack_0 <= ackL_unguarded(3);
      LOAD_pad_2216_load_0_ack_0 <= ackL_unguarded(2);
      LOAD_pad_2627_load_0_ack_0 <= ackL_unguarded(1);
      LOAD_pad_3030_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= LOAD_pad_1000_load_0_req_1;
      reqR_unguarded(6) <= LOAD_pad_512_load_0_req_1;
      reqR_unguarded(5) <= LOAD_pad_3441_load_0_req_1;
      reqR_unguarded(4) <= LOAD_pad_1408_load_0_req_1;
      reqR_unguarded(3) <= LOAD_pad_1813_load_0_req_1;
      reqR_unguarded(2) <= LOAD_pad_2216_load_0_req_1;
      reqR_unguarded(1) <= LOAD_pad_2627_load_0_req_1;
      reqR_unguarded(0) <= LOAD_pad_3030_load_0_req_1;
      LOAD_pad_1000_load_0_ack_1 <= ackR_unguarded(7);
      LOAD_pad_512_load_0_ack_1 <= ackR_unguarded(6);
      LOAD_pad_3441_load_0_ack_1 <= ackR_unguarded(5);
      LOAD_pad_1408_load_0_ack_1 <= ackR_unguarded(4);
      LOAD_pad_1813_load_0_ack_1 <= ackR_unguarded(3);
      LOAD_pad_2216_load_0_ack_1 <= ackR_unguarded(2);
      LOAD_pad_2627_load_0_ack_1 <= ackR_unguarded(1);
      LOAD_pad_3030_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_pad_1000_word_address_0 & LOAD_pad_512_word_address_0 & LOAD_pad_3441_word_address_0 & LOAD_pad_1408_word_address_0 & LOAD_pad_1813_word_address_0 & LOAD_pad_2216_word_address_0 & LOAD_pad_2627_word_address_0 & LOAD_pad_3030_word_address_0;
      LOAD_pad_1000_data_0 <= data_out(63 downto 56);
      LOAD_pad_512_data_0 <= data_out(55 downto 48);
      LOAD_pad_3441_data_0 <= data_out(47 downto 40);
      LOAD_pad_1408_data_0 <= data_out(39 downto 32);
      LOAD_pad_1813_data_0 <= data_out(31 downto 24);
      LOAD_pad_2216_data_0 <= data_out(23 downto 16);
      LOAD_pad_2627_data_0 <= data_out(15 downto 8);
      LOAD_pad_3030_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(0 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(7 downto 0),
          mtag => memory_space_3_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_856_load_0 ptr_deref_1265_load_0 ptr_deref_3295_load_0 ptr_deref_1679_load_0 ptr_deref_2077_load_0 ptr_deref_2493_load_0 ptr_deref_2891_load_0 ptr_deref_3705_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(111 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      reqL_unguarded(7) <= ptr_deref_856_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_1265_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_3295_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1679_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_2077_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_2493_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2891_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3705_load_0_req_0;
      ptr_deref_856_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_1265_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_3295_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1679_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_2077_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_2493_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2891_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3705_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_856_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_1265_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_3295_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1679_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_2077_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_2493_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2891_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3705_load_0_req_1;
      ptr_deref_856_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_1265_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_3295_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1679_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_2077_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_2493_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2891_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3705_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_856_word_address_0 & ptr_deref_1265_word_address_0 & ptr_deref_3295_word_address_0 & ptr_deref_1679_word_address_0 & ptr_deref_2077_word_address_0 & ptr_deref_2493_word_address_0 & ptr_deref_2891_word_address_0 & ptr_deref_3705_word_address_0;
      ptr_deref_856_data_0 <= data_out(511 downto 448);
      ptr_deref_1265_data_0 <= data_out(447 downto 384);
      ptr_deref_3295_data_0 <= data_out(383 downto 320);
      ptr_deref_1679_data_0 <= data_out(319 downto 256);
      ptr_deref_2077_data_0 <= data_out(255 downto 192);
      ptr_deref_2493_data_0 <= data_out(191 downto 128);
      ptr_deref_2891_data_0 <= data_out(127 downto 64);
      ptr_deref_3705_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : STORE_pad_242_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_pad_242_store_0_req_0;
      STORE_pad_242_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_pad_242_store_0_req_1;
      STORE_pad_242_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_pad_242_word_address_0;
      data_in <= STORE_pad_242_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(0 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_772_store_0 ptr_deref_1181_store_0 ptr_deref_880_store_0 ptr_deref_1289_store_0 ptr_deref_3211_store_0 ptr_deref_3319_store_0 ptr_deref_1595_store_0 ptr_deref_1703_store_0 ptr_deref_1993_store_0 ptr_deref_2101_store_0 ptr_deref_2409_store_0 ptr_deref_2517_store_0 ptr_deref_2807_store_0 ptr_deref_2915_store_0 ptr_deref_3621_store_0 ptr_deref_3729_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(223 downto 0);
      signal data_in: std_logic_vector(1023 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 15 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(15 downto 0) := (15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      reqL_unguarded(15) <= ptr_deref_772_store_0_req_0;
      reqL_unguarded(14) <= ptr_deref_1181_store_0_req_0;
      reqL_unguarded(13) <= ptr_deref_880_store_0_req_0;
      reqL_unguarded(12) <= ptr_deref_1289_store_0_req_0;
      reqL_unguarded(11) <= ptr_deref_3211_store_0_req_0;
      reqL_unguarded(10) <= ptr_deref_3319_store_0_req_0;
      reqL_unguarded(9) <= ptr_deref_1595_store_0_req_0;
      reqL_unguarded(8) <= ptr_deref_1703_store_0_req_0;
      reqL_unguarded(7) <= ptr_deref_1993_store_0_req_0;
      reqL_unguarded(6) <= ptr_deref_2101_store_0_req_0;
      reqL_unguarded(5) <= ptr_deref_2409_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_2517_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_2807_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_2915_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_3621_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3729_store_0_req_0;
      ptr_deref_772_store_0_ack_0 <= ackL_unguarded(15);
      ptr_deref_1181_store_0_ack_0 <= ackL_unguarded(14);
      ptr_deref_880_store_0_ack_0 <= ackL_unguarded(13);
      ptr_deref_1289_store_0_ack_0 <= ackL_unguarded(12);
      ptr_deref_3211_store_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_3319_store_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_1595_store_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_1703_store_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_1993_store_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_2101_store_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_2409_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_2517_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_2807_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_2915_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_3621_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3729_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(15) <= ptr_deref_772_store_0_req_1;
      reqR_unguarded(14) <= ptr_deref_1181_store_0_req_1;
      reqR_unguarded(13) <= ptr_deref_880_store_0_req_1;
      reqR_unguarded(12) <= ptr_deref_1289_store_0_req_1;
      reqR_unguarded(11) <= ptr_deref_3211_store_0_req_1;
      reqR_unguarded(10) <= ptr_deref_3319_store_0_req_1;
      reqR_unguarded(9) <= ptr_deref_1595_store_0_req_1;
      reqR_unguarded(8) <= ptr_deref_1703_store_0_req_1;
      reqR_unguarded(7) <= ptr_deref_1993_store_0_req_1;
      reqR_unguarded(6) <= ptr_deref_2101_store_0_req_1;
      reqR_unguarded(5) <= ptr_deref_2409_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_2517_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_2807_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_2915_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_3621_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3729_store_0_req_1;
      ptr_deref_772_store_0_ack_1 <= ackR_unguarded(15);
      ptr_deref_1181_store_0_ack_1 <= ackR_unguarded(14);
      ptr_deref_880_store_0_ack_1 <= ackR_unguarded(13);
      ptr_deref_1289_store_0_ack_1 <= ackR_unguarded(12);
      ptr_deref_3211_store_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_3319_store_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_1595_store_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_1703_store_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_1993_store_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_2101_store_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_2409_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_2517_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_2807_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_2915_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_3621_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3729_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_6: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_6", num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_7: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_7", num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_8: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_8", num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_9: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_9", num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_10: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_10", num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_11: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_11", num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_12: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_12", num_slots => 1) -- 
        port map (req => reqL_unregulated(12), -- 
          ack => ackL_unregulated(12),
          regulated_req => reqL(12),
          regulated_ack => ackL(12),
          release_req => reqR(12),
          release_ack => ackR(12),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_13: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_13", num_slots => 1) -- 
        port map (req => reqL_unregulated(13), -- 
          ack => ackL_unregulated(13),
          regulated_req => reqL(13),
          regulated_ack => ackL(13),
          release_req => reqR(13),
          release_ack => ackR(13),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_14: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_14", num_slots => 1) -- 
        port map (req => reqL_unregulated(14), -- 
          ack => ackL_unregulated(14),
          regulated_req => reqL(14),
          regulated_ack => ackL(14),
          release_req => reqR(14),
          release_ack => ackR(14),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_15: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_15", num_slots => 1) -- 
        port map (req => reqL_unregulated(15), -- 
          ack => ackL_unregulated(15),
          regulated_req => reqL(15),
          regulated_ack => ackL(15),
          release_req => reqR(15),
          release_ack => ackR(15),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_772_word_address_0 & ptr_deref_1181_word_address_0 & ptr_deref_880_word_address_0 & ptr_deref_1289_word_address_0 & ptr_deref_3211_word_address_0 & ptr_deref_3319_word_address_0 & ptr_deref_1595_word_address_0 & ptr_deref_1703_word_address_0 & ptr_deref_1993_word_address_0 & ptr_deref_2101_word_address_0 & ptr_deref_2409_word_address_0 & ptr_deref_2517_word_address_0 & ptr_deref_2807_word_address_0 & ptr_deref_2915_word_address_0 & ptr_deref_3621_word_address_0 & ptr_deref_3729_word_address_0;
      data_in <= ptr_deref_772_data_0 & ptr_deref_1181_data_0 & ptr_deref_880_data_0 & ptr_deref_1289_data_0 & ptr_deref_3211_data_0 & ptr_deref_3319_data_0 & ptr_deref_1595_data_0 & ptr_deref_1703_data_0 & ptr_deref_1993_data_0 & ptr_deref_2101_data_0 & ptr_deref_2409_data_0 & ptr_deref_2517_data_0 & ptr_deref_2807_data_0 & ptr_deref_2915_data_0 & ptr_deref_3621_data_0 & ptr_deref_3729_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(21 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 16,
          detailed_buffering_per_output => outBUFs,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_487_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_487_store_0_req_0;
      ptr_deref_487_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_487_store_0_req_1;
      ptr_deref_487_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_487_word_address_0;
      data_in <= ptr_deref_487_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_zeropad_input_pipe_237_inst RPIPE_zeropad_input_pipe_240_inst RPIPE_zeropad_input_pipe_367_inst RPIPE_zeropad_input_pipe_234_inst RPIPE_zeropad_input_pipe_252_inst RPIPE_zeropad_input_pipe_231_inst RPIPE_zeropad_input_pipe_228_inst RPIPE_zeropad_input_pipe_225_inst RPIPE_zeropad_input_pipe_354_inst RPIPE_zeropad_input_pipe_249_inst RPIPE_zeropad_input_pipe_246_inst RPIPE_zeropad_input_pipe_385_inst RPIPE_zeropad_input_pipe_403_inst RPIPE_zeropad_input_pipe_421_inst RPIPE_zeropad_input_pipe_439_inst RPIPE_zeropad_input_pipe_457_inst RPIPE_zeropad_input_pipe_475_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(135 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 16 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 16 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 16 downto 0);
      signal guard_vector : std_logic_vector( 16 downto 0);
      constant outBUFs : IntegerArray(16 downto 0) := (16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(16 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false);
      constant guardBuffering: IntegerArray(16 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2);
      -- 
    begin -- 
      reqL_unguarded(16) <= RPIPE_zeropad_input_pipe_237_inst_req_0;
      reqL_unguarded(15) <= RPIPE_zeropad_input_pipe_240_inst_req_0;
      reqL_unguarded(14) <= RPIPE_zeropad_input_pipe_367_inst_req_0;
      reqL_unguarded(13) <= RPIPE_zeropad_input_pipe_234_inst_req_0;
      reqL_unguarded(12) <= RPIPE_zeropad_input_pipe_252_inst_req_0;
      reqL_unguarded(11) <= RPIPE_zeropad_input_pipe_231_inst_req_0;
      reqL_unguarded(10) <= RPIPE_zeropad_input_pipe_228_inst_req_0;
      reqL_unguarded(9) <= RPIPE_zeropad_input_pipe_225_inst_req_0;
      reqL_unguarded(8) <= RPIPE_zeropad_input_pipe_354_inst_req_0;
      reqL_unguarded(7) <= RPIPE_zeropad_input_pipe_249_inst_req_0;
      reqL_unguarded(6) <= RPIPE_zeropad_input_pipe_246_inst_req_0;
      reqL_unguarded(5) <= RPIPE_zeropad_input_pipe_385_inst_req_0;
      reqL_unguarded(4) <= RPIPE_zeropad_input_pipe_403_inst_req_0;
      reqL_unguarded(3) <= RPIPE_zeropad_input_pipe_421_inst_req_0;
      reqL_unguarded(2) <= RPIPE_zeropad_input_pipe_439_inst_req_0;
      reqL_unguarded(1) <= RPIPE_zeropad_input_pipe_457_inst_req_0;
      reqL_unguarded(0) <= RPIPE_zeropad_input_pipe_475_inst_req_0;
      RPIPE_zeropad_input_pipe_237_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_zeropad_input_pipe_240_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_zeropad_input_pipe_367_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_zeropad_input_pipe_234_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_zeropad_input_pipe_252_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_zeropad_input_pipe_231_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_zeropad_input_pipe_228_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_zeropad_input_pipe_225_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_zeropad_input_pipe_354_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_zeropad_input_pipe_249_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_zeropad_input_pipe_246_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_zeropad_input_pipe_385_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_zeropad_input_pipe_403_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_zeropad_input_pipe_421_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_zeropad_input_pipe_439_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_zeropad_input_pipe_457_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_zeropad_input_pipe_475_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(16) <= RPIPE_zeropad_input_pipe_237_inst_req_1;
      reqR_unguarded(15) <= RPIPE_zeropad_input_pipe_240_inst_req_1;
      reqR_unguarded(14) <= RPIPE_zeropad_input_pipe_367_inst_req_1;
      reqR_unguarded(13) <= RPIPE_zeropad_input_pipe_234_inst_req_1;
      reqR_unguarded(12) <= RPIPE_zeropad_input_pipe_252_inst_req_1;
      reqR_unguarded(11) <= RPIPE_zeropad_input_pipe_231_inst_req_1;
      reqR_unguarded(10) <= RPIPE_zeropad_input_pipe_228_inst_req_1;
      reqR_unguarded(9) <= RPIPE_zeropad_input_pipe_225_inst_req_1;
      reqR_unguarded(8) <= RPIPE_zeropad_input_pipe_354_inst_req_1;
      reqR_unguarded(7) <= RPIPE_zeropad_input_pipe_249_inst_req_1;
      reqR_unguarded(6) <= RPIPE_zeropad_input_pipe_246_inst_req_1;
      reqR_unguarded(5) <= RPIPE_zeropad_input_pipe_385_inst_req_1;
      reqR_unguarded(4) <= RPIPE_zeropad_input_pipe_403_inst_req_1;
      reqR_unguarded(3) <= RPIPE_zeropad_input_pipe_421_inst_req_1;
      reqR_unguarded(2) <= RPIPE_zeropad_input_pipe_439_inst_req_1;
      reqR_unguarded(1) <= RPIPE_zeropad_input_pipe_457_inst_req_1;
      reqR_unguarded(0) <= RPIPE_zeropad_input_pipe_475_inst_req_1;
      RPIPE_zeropad_input_pipe_237_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_zeropad_input_pipe_240_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_zeropad_input_pipe_367_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_zeropad_input_pipe_234_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_zeropad_input_pipe_252_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_zeropad_input_pipe_231_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_zeropad_input_pipe_228_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_zeropad_input_pipe_225_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_zeropad_input_pipe_354_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_zeropad_input_pipe_249_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_zeropad_input_pipe_246_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_zeropad_input_pipe_385_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_zeropad_input_pipe_403_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_zeropad_input_pipe_421_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_zeropad_input_pipe_439_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_zeropad_input_pipe_457_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_zeropad_input_pipe_475_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      call4_238 <= data_out(135 downto 128);
      call5_241 <= data_out(127 downto 120);
      call23_368 <= data_out(119 downto 112);
      call3_235 <= data_out(111 downto 104);
      call8_253 <= data_out(103 downto 96);
      call2_232 <= data_out(95 downto 88);
      call1_229 <= data_out(87 downto 80);
      call_226 <= data_out(79 downto 72);
      call20_355 <= data_out(71 downto 64);
      call7_250 <= data_out(63 downto 56);
      call6_247 <= data_out(55 downto 48);
      call28_386 <= data_out(47 downto 40);
      call34_404 <= data_out(39 downto 32);
      call40_422 <= data_out(31 downto 24);
      call46_440 <= data_out(23 downto 16);
      call52_458 <= data_out(15 downto 8);
      call58_476 <= data_out(7 downto 0);
      zeropad_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "zeropad_input_pipe_read_0_gI", nreqs => 17, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      zeropad_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "zeropad_input_pipe_read_0", data_width => 8,  num_reqs => 17,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => zeropad_input_pipe_pipe_read_req(0),
          oack => zeropad_input_pipe_pipe_read_ack(0),
          odata => zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_3857_call 
    sendOutput_call_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_3857_call_req_0;
      call_stmt_3857_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_3857_call_req_1;
      call_stmt_3857_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_0_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul1794_3855;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          dataR => sendOutput_call_data(31 downto 0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(21 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(21 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_2
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(4 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_size :  std_logic_vector(31 downto 0);
  signal sendOutput_in_args    : std_logic_vector(31 downto 0);
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_data: std_logic_vector(31 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module zeropad3D
  component zeropad3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(21 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(3 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_data : out  std_logic_vector(31 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D
  signal zeropad3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_start_req : std_logic;
  signal zeropad3D_start_ack : std_logic;
  signal zeropad3D_fin_req   : std_logic;
  signal zeropad3D_fin_ack : std_logic;
  -- aggregate signals for read from pipe zeropad_input_pipe
  signal zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe zeropad_output_pipe
  signal zeropad_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal zeropad_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal zeropad_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module sendOutput
  sendOutput_size <= sendOutput_in_args(31 downto 0);
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_data  => sendOutput_call_data,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      call_mdata => sendOutput_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendOutput_size,
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(21 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(4 downto 0),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(0 downto 0),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(0 downto 0),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module zeropad3D
  zeropad3D_instance:zeropad3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_start_req,
      start_ack => zeropad3D_start_ack,
      fin_req => zeropad3D_fin_req,
      fin_ack => zeropad3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(0 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(20 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(7 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(3 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(21 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(4 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(3 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(0 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(7 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(20 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 0),
      zeropad_input_pipe_pipe_read_req => zeropad_input_pipe_pipe_read_req(0 downto 0),
      zeropad_input_pipe_pipe_read_ack => zeropad_input_pipe_pipe_read_ack(0 downto 0),
      zeropad_input_pipe_pipe_read_data => zeropad_input_pipe_pipe_read_data(7 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_data => sendOutput_call_data(31 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      tag_in => zeropad3D_tag_in,
      tag_out => zeropad3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_tag_in <= (others => '0');
  zeropad3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_start_req, start_ack => zeropad3D_start_ack,  fin_req => zeropad3D_fin_req,  fin_ack => zeropad3D_fin_ack);
  zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_input_pipe_pipe_read_req,
      read_ack => zeropad_input_pipe_pipe_read_ack,
      read_data => zeropad_input_pipe_pipe_read_data,
      write_req => zeropad_input_pipe_pipe_write_req,
      write_ack => zeropad_input_pipe_pipe_write_ack,
      write_data => zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_output_pipe_pipe_read_req,
      read_ack => zeropad_output_pipe_pipe_read_ack,
      read_data => zeropad_output_pipe_pipe_read_data,
      write_req => zeropad_output_pipe_pipe_write_req,
      write_ack => zeropad_output_pipe_pipe_write_ack,
      write_data => zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 5,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
